--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_73986f767e994888.vhd when simulating
-- the core, addsb_11_0_73986f767e994888. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_73986f767e994888 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END addsb_11_0_73986f767e994888;

ARCHITECTURE addsb_11_0_73986f767e994888_a OF addsb_11_0_73986f767e994888 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_73986f767e994888
  PORT (
    a : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_73986f767e994888 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 10,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "0000000000",
      c_b_width => 10,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 10,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_73986f767e994888
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_73986f767e994888_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_8dc9188fad4d9a9c.vhd when simulating
-- the core, addsb_11_0_8dc9188fad4d9a9c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_8dc9188fad4d9a9c IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END addsb_11_0_8dc9188fad4d9a9c;

ARCHITECTURE addsb_11_0_8dc9188fad4d9a9c_a OF addsb_11_0_8dc9188fad4d9a9c IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_8dc9188fad4d9a9c
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_8dc9188fad4d9a9c USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 9,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "000000000",
      c_b_width => 9,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 9,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_8dc9188fad4d9a9c
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_8dc9188fad4d9a9c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_913f4bce6842c815.vhd when simulating
-- the core, addsb_11_0_913f4bce6842c815. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_913f4bce6842c815 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END addsb_11_0_913f4bce6842c815;

ARCHITECTURE addsb_11_0_913f4bce6842c815_a OF addsb_11_0_913f4bce6842c815 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_913f4bce6842c815
  PORT (
    a : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(12 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_913f4bce6842c815 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 13,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "0000000000000",
      c_b_width => 13,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 13,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_913f4bce6842c815
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_913f4bce6842c815_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_a52ead9b8a3c1e76.vhd when simulating
-- the core, addsb_11_0_a52ead9b8a3c1e76. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_a52ead9b8a3c1e76 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END addsb_11_0_a52ead9b8a3c1e76;

ARCHITECTURE addsb_11_0_a52ead9b8a3c1e76_a OF addsb_11_0_a52ead9b8a3c1e76 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_a52ead9b8a3c1e76
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_a52ead9b8a3c1e76 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 9,
      c_add_mode => 1,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 0,
      c_b_value => "000000000",
      c_b_width => 9,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 9,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_a52ead9b8a3c1e76
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_a52ead9b8a3c1e76_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file axififo_fg92_4d50ffea04713b7c.vhd when simulating
-- the core, axififo_fg92_4d50ffea04713b7c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY axififo_fg92_4d50ffea04713b7c IS
  PORT (
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    s_axis_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    m_axis_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
  );
END axififo_fg92_4d50ffea04713b7c;

ARCHITECTURE axififo_fg92_4d50ffea04713b7c_a OF axififo_fg92_4d50ffea04713b7c IS
-- synthesis translate_off
COMPONENT wrapped_axififo_fg92_4d50ffea04713b7c
  PORT (
    s_aclk : IN STD_LOGIC;
    s_aresetn : IN STD_LOGIC;
    s_axis_tvalid : IN STD_LOGIC;
    s_axis_tready : OUT STD_LOGIC;
    s_axis_tdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    s_axis_tlast : IN STD_LOGIC;
    s_axis_tuser : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    m_axis_tvalid : OUT STD_LOGIC;
    m_axis_tready : IN STD_LOGIC;
    m_axis_tdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    m_axis_tlast : OUT STD_LOGIC;
    m_axis_tuser : OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_axififo_fg92_4d50ffea04713b7c USE ENTITY XilinxCoreLib.fifo_generator_v9_3(behavioral)
    GENERIC MAP (
      c_add_ngc_constraint => 0,
      c_application_type_axis => 0,
      c_application_type_rach => 0,
      c_application_type_rdch => 0,
      c_application_type_wach => 0,
      c_application_type_wdch => 0,
      c_application_type_wrch => 0,
      c_axi_addr_width => 32,
      c_axi_aruser_width => 1,
      c_axi_awuser_width => 1,
      c_axi_buser_width => 1,
      c_axi_data_width => 64,
      c_axi_id_width => 4,
      c_axi_ruser_width => 1,
      c_axi_type => 0,
      c_axi_wuser_width => 1,
      c_axis_tdata_width => 32,
      c_axis_tdest_width => 4,
      c_axis_tid_width => 8,
      c_axis_tkeep_width => 4,
      c_axis_tstrb_width => 4,
      c_axis_tuser_width => 1,
      c_axis_type => 0,
      c_common_clock => 1,
      c_count_type => 0,
      c_data_count_width => 10,
      c_default_value => "BlankString",
      c_din_width => 18,
      c_din_width_axis => 34,
      c_din_width_rach => 32,
      c_din_width_rdch => 64,
      c_din_width_wach => 32,
      c_din_width_wdch => 64,
      c_din_width_wrch => 2,
      c_dout_rst_val => "0",
      c_dout_width => 18,
      c_enable_rlocs => 0,
      c_enable_rst_sync => 1,
      c_error_injection_type => 0,
      c_error_injection_type_axis => 0,
      c_error_injection_type_rach => 0,
      c_error_injection_type_rdch => 0,
      c_error_injection_type_wach => 0,
      c_error_injection_type_wdch => 0,
      c_error_injection_type_wrch => 0,
      c_family => "virtex6",
      c_full_flags_rst_val => 1,
      c_has_almost_empty => 0,
      c_has_almost_full => 0,
      c_has_axi_aruser => 0,
      c_has_axi_awuser => 0,
      c_has_axi_buser => 0,
      c_has_axi_rd_channel => 0,
      c_has_axi_ruser => 0,
      c_has_axi_wr_channel => 0,
      c_has_axi_wuser => 0,
      c_has_axis_tdata => 1,
      c_has_axis_tdest => 0,
      c_has_axis_tid => 0,
      c_has_axis_tkeep => 0,
      c_has_axis_tlast => 1,
      c_has_axis_tready => 1,
      c_has_axis_tstrb => 0,
      c_has_axis_tuser => 1,
      c_has_backup => 0,
      c_has_data_count => 0,
      c_has_data_counts_axis => 0,
      c_has_data_counts_rach => 0,
      c_has_data_counts_rdch => 0,
      c_has_data_counts_wach => 0,
      c_has_data_counts_wdch => 0,
      c_has_data_counts_wrch => 0,
      c_has_int_clk => 0,
      c_has_master_ce => 0,
      c_has_meminit_file => 0,
      c_has_overflow => 0,
      c_has_prog_flags_axis => 0,
      c_has_prog_flags_rach => 0,
      c_has_prog_flags_rdch => 0,
      c_has_prog_flags_wach => 0,
      c_has_prog_flags_wdch => 0,
      c_has_prog_flags_wrch => 0,
      c_has_rd_data_count => 0,
      c_has_rd_rst => 0,
      c_has_rst => 1,
      c_has_slave_ce => 0,
      c_has_srst => 0,
      c_has_underflow => 0,
      c_has_valid => 0,
      c_has_wr_ack => 0,
      c_has_wr_data_count => 0,
      c_has_wr_rst => 0,
      c_implementation_type => 0,
      c_implementation_type_axis => 1,
      c_implementation_type_rach => 2,
      c_implementation_type_rdch => 1,
      c_implementation_type_wach => 2,
      c_implementation_type_wdch => 1,
      c_implementation_type_wrch => 2,
      c_init_wr_pntr_val => 0,
      c_interface_type => 1,
      c_memory_type => 1,
      c_mif_file_name => "BlankString",
      c_msgon_val => 1,
      c_optimization_mode => 0,
      c_overflow_low => 0,
      c_preload_latency => 1,
      c_preload_regs => 0,
      c_prim_fifo_type => "4kx4",
      c_prog_empty_thresh_assert_val => 2,
      c_prog_empty_thresh_assert_val_axis => 62,
      c_prog_empty_thresh_assert_val_rach => 14,
      c_prog_empty_thresh_assert_val_rdch => 1022,
      c_prog_empty_thresh_assert_val_wach => 14,
      c_prog_empty_thresh_assert_val_wdch => 1022,
      c_prog_empty_thresh_assert_val_wrch => 14,
      c_prog_empty_thresh_negate_val => 3,
      c_prog_empty_type => 0,
      c_prog_empty_type_axis => 0,
      c_prog_empty_type_rach => 0,
      c_prog_empty_type_rdch => 0,
      c_prog_empty_type_wach => 0,
      c_prog_empty_type_wdch => 0,
      c_prog_empty_type_wrch => 0,
      c_prog_full_thresh_assert_val => 1022,
      c_prog_full_thresh_assert_val_axis => 63,
      c_prog_full_thresh_assert_val_rach => 15,
      c_prog_full_thresh_assert_val_rdch => 1023,
      c_prog_full_thresh_assert_val_wach => 15,
      c_prog_full_thresh_assert_val_wdch => 1023,
      c_prog_full_thresh_assert_val_wrch => 15,
      c_prog_full_thresh_negate_val => 1021,
      c_prog_full_type => 0,
      c_prog_full_type_axis => 0,
      c_prog_full_type_rach => 0,
      c_prog_full_type_rdch => 0,
      c_prog_full_type_wach => 0,
      c_prog_full_type_wdch => 0,
      c_prog_full_type_wrch => 0,
      c_rach_type => 0,
      c_rd_data_count_width => 10,
      c_rd_depth => 1024,
      c_rd_freq => 1,
      c_rd_pntr_width => 10,
      c_rdch_type => 0,
      c_reg_slice_mode_axis => 0,
      c_reg_slice_mode_rach => 0,
      c_reg_slice_mode_rdch => 0,
      c_reg_slice_mode_wach => 0,
      c_reg_slice_mode_wdch => 0,
      c_reg_slice_mode_wrch => 0,
      c_synchronizer_stage => 2,
      c_underflow_low => 0,
      c_use_common_overflow => 0,
      c_use_common_underflow => 0,
      c_use_default_settings => 0,
      c_use_dout_rst => 1,
      c_use_ecc => 0,
      c_use_ecc_axis => 0,
      c_use_ecc_rach => 0,
      c_use_ecc_rdch => 0,
      c_use_ecc_wach => 0,
      c_use_ecc_wdch => 0,
      c_use_ecc_wrch => 0,
      c_use_embedded_reg => 0,
      c_use_fifo16_flags => 0,
      c_use_fwft_data_count => 0,
      c_valid_low => 0,
      c_wach_type => 0,
      c_wdch_type => 0,
      c_wr_ack_low => 0,
      c_wr_data_count_width => 10,
      c_wr_depth => 1024,
      c_wr_depth_axis => 64,
      c_wr_depth_rach => 16,
      c_wr_depth_rdch => 1024,
      c_wr_depth_wach => 16,
      c_wr_depth_wdch => 1024,
      c_wr_depth_wrch => 16,
      c_wr_freq => 1,
      c_wr_pntr_width => 10,
      c_wr_pntr_width_axis => 6,
      c_wr_pntr_width_rach => 4,
      c_wr_pntr_width_rdch => 10,
      c_wr_pntr_width_wach => 4,
      c_wr_pntr_width_wdch => 10,
      c_wr_pntr_width_wrch => 4,
      c_wr_response_latency => 1,
      c_wrch_type => 0
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_axififo_fg92_4d50ffea04713b7c
  PORT MAP (
    s_aclk => s_aclk,
    s_aresetn => s_aresetn,
    s_axis_tvalid => s_axis_tvalid,
    s_axis_tready => s_axis_tready,
    s_axis_tdata => s_axis_tdata,
    s_axis_tlast => s_axis_tlast,
    s_axis_tuser => s_axis_tuser,
    m_axis_tvalid => m_axis_tvalid,
    m_axis_tready => m_axis_tready,
    m_axis_tdata => m_axis_tdata,
    m_axis_tlast => m_axis_tlast,
    m_axis_tuser => m_axis_tuser
  );
-- synthesis translate_on

END axififo_fg92_4d50ffea04713b7c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_28f68c2bb9b4d938.vhd when simulating
-- the core, bmg_72_28f68c2bb9b4d938. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_28f68c2bb9b4d938 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END bmg_72_28f68c2bb9b4d938;

ARCHITECTURE bmg_72_28f68c2bb9b4d938_a OF bmg_72_28f68c2bb9b4d938 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_28f68c2bb9b4d938
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_28f68c2bb9b4d938 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 8,
      c_addrb_width => 8,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_28f68c2bb9b4d938.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 192,
      c_read_depth_b => 192,
      c_read_width_a => 8,
      c_read_width_b => 8,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 192,
      c_write_depth_b => 192,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 8,
      c_write_width_b => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_28f68c2bb9b4d938
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_28f68c2bb9b4d938_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_324b883165919716.vhd when simulating
-- the core, bmg_72_324b883165919716. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_324b883165919716 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END bmg_72_324b883165919716;

ARCHITECTURE bmg_72_324b883165919716_a OF bmg_72_324b883165919716 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_324b883165919716
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_324b883165919716 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 9,
      c_addrb_width => 9,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_324b883165919716.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 288,
      c_read_depth_b => 288,
      c_read_width_a => 9,
      c_read_width_b => 9,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 288,
      c_write_depth_b => 288,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 9,
      c_write_width_b => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_324b883165919716
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_324b883165919716_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_3628803596b5ca22.vhd when simulating
-- the core, bmg_72_3628803596b5ca22. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_3628803596b5ca22 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END bmg_72_3628803596b5ca22;

ARCHITECTURE bmg_72_3628803596b5ca22_a OF bmg_72_3628803596b5ca22 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_3628803596b5ca22
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_3628803596b5ca22 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 7,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_3628803596b5ca22.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 96,
      c_read_depth_b => 96,
      c_read_width_a => 7,
      c_read_width_b => 7,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 96,
      c_write_depth_b => 96,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 7,
      c_write_width_b => 7,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_3628803596b5ca22
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_3628803596b5ca22_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_376dc060ca4075f2.vhd when simulating
-- the core, bmg_72_376dc060ca4075f2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_376dc060ca4075f2 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END bmg_72_376dc060ca4075f2;

ARCHITECTURE bmg_72_376dc060ca4075f2_a OF bmg_72_376dc060ca4075f2 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_376dc060ca4075f2
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_376dc060ca4075f2 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 8,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_376dc060ca4075f2.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 256,
      c_read_depth_b => 128,
      c_read_width_a => 1,
      c_read_width_b => 2,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 256,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 1,
      c_write_width_b => 2,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_376dc060ca4075f2
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_376dc060ca4075f2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_41985f385eaacb3e.vhd when simulating
-- the core, bmg_72_41985f385eaacb3e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_41985f385eaacb3e IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
  );
END bmg_72_41985f385eaacb3e;

ARCHITECTURE bmg_72_41985f385eaacb3e_a OF bmg_72_41985f385eaacb3e IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_41985f385eaacb3e
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_41985f385eaacb3e USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 7,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_41985f385eaacb3e.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 128,
      c_read_depth_b => 128,
      c_read_width_a => 1,
      c_read_width_b => 1,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 128,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 1,
      c_write_width_b => 1,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_41985f385eaacb3e
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_41985f385eaacb3e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_7ec9033b751d2879.vhd when simulating
-- the core, bmg_72_7ec9033b751d2879. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_7ec9033b751d2879 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END bmg_72_7ec9033b751d2879;

ARCHITECTURE bmg_72_7ec9033b751d2879_a OF bmg_72_7ec9033b751d2879 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_7ec9033b751d2879
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_7ec9033b751d2879 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 9,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_7ec9033b751d2879.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 512,
      c_read_depth_b => 128,
      c_read_width_a => 1,
      c_read_width_b => 4,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 512,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 1,
      c_write_width_b => 4,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_7ec9033b751d2879
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_7ec9033b751d2879_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_da153342fc52049b.vhd when simulating
-- the core, bmg_72_da153342fc52049b. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_da153342fc52049b IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END bmg_72_da153342fc52049b;

ARCHITECTURE bmg_72_da153342fc52049b_a OF bmg_72_da153342fc52049b IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_da153342fc52049b
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    clkb : IN STD_LOGIC;
    enb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_da153342fc52049b USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 10,
      c_addrb_width => 7,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 1,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 1,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_da153342fc52049b.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 2,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 1024,
      c_read_depth_b => 128,
      c_read_width_a => 1,
      c_read_width_b => 8,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 1024,
      c_write_depth_b => 128,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 1,
      c_write_width_b => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_da153342fc52049b
  PORT MAP (
    clka => clka,
    ena => ena,
    wea => wea,
    addra => addra,
    dina => dina,
    douta => douta,
    clkb => clkb,
    enb => enb,
    web => web,
    addrb => addrb,
    dinb => dinb,
    doutb => doutb
  );
-- synthesis translate_on

END bmg_72_da153342fc52049b_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file bmg_72_f580ae3be5511d30.vhd when simulating
-- the core, bmg_72_f580ae3be5511d30. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY bmg_72_f580ae3be5511d30 IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END bmg_72_f580ae3be5511d30;

ARCHITECTURE bmg_72_f580ae3be5511d30_a OF bmg_72_f580ae3be5511d30 IS
-- synthesis translate_off
COMPONENT wrapped_bmg_72_f580ae3be5511d30
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_bmg_72_f580ae3be5511d30 USE ENTITY XilinxCoreLib.blk_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addra_width => 6,
      c_addrb_width => 6,
      c_algorithm => 1,
      c_axi_id_width => 4,
      c_axi_slave_type => 0,
      c_axi_type => 1,
      c_byte_size => 9,
      c_common_clk => 0,
      c_default_data => "0",
      c_disable_warn_bhv_coll => 0,
      c_disable_warn_bhv_range => 0,
      c_enable_32bit_address => 0,
      c_family => "virtex6",
      c_has_axi_id => 0,
      c_has_ena => 1,
      c_has_enb => 0,
      c_has_injecterr => 0,
      c_has_mem_output_regs_a => 0,
      c_has_mem_output_regs_b => 0,
      c_has_mux_output_regs_a => 0,
      c_has_mux_output_regs_b => 0,
      c_has_regcea => 0,
      c_has_regceb => 0,
      c_has_rsta => 0,
      c_has_rstb => 0,
      c_has_softecc_input_regs_a => 0,
      c_has_softecc_output_regs_b => 0,
      c_init_file_name => "bmg_72_f580ae3be5511d30.mif",
      c_inita_val => "0",
      c_initb_val => "0",
      c_interface_type => 0,
      c_load_init_file => 1,
      c_mem_type => 3,
      c_mux_pipeline_stages => 0,
      c_prim_type => 1,
      c_read_depth_a => 48,
      c_read_depth_b => 48,
      c_read_width_a => 6,
      c_read_width_b => 6,
      c_rst_priority_a => "CE",
      c_rst_priority_b => "CE",
      c_rst_type => "SYNC",
      c_rstram_a => 0,
      c_rstram_b => 0,
      c_sim_collision_check => "ALL",
      c_use_byte_wea => 0,
      c_use_byte_web => 0,
      c_use_default_data => 0,
      c_use_ecc => 0,
      c_use_softecc => 0,
      c_wea_width => 1,
      c_web_width => 1,
      c_write_depth_a => 48,
      c_write_depth_b => 48,
      c_write_mode_a => "WRITE_FIRST",
      c_write_mode_b => "WRITE_FIRST",
      c_write_width_a => 6,
      c_write_width_b => 6,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_bmg_72_f580ae3be5511d30
  PORT MAP (
    clka => clka,
    ena => ena,
    addra => addra,
    douta => douta
  );
-- synthesis translate_on

END bmg_72_f580ae3be5511d30_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_36e2bb554c95560d.vhd when simulating
-- the core, cntr_11_0_36e2bb554c95560d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_36e2bb554c95560d IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END cntr_11_0_36e2bb554c95560d;

ARCHITECTURE cntr_11_0_36e2bb554c95560d_a OF cntr_11_0_36e2bb554c95560d IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_36e2bb554c95560d
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_36e2bb554c95560d USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_36e2bb554c95560d
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_36e2bb554c95560d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_6454489cfe866515.vhd when simulating
-- the core, cntr_11_0_6454489cfe866515. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_6454489cfe866515 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END cntr_11_0_6454489cfe866515;

ARCHITECTURE cntr_11_0_6454489cfe866515_a OF cntr_11_0_6454489cfe866515 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_6454489cfe866515
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_6454489cfe866515 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 2,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_6454489cfe866515
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_6454489cfe866515_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_86806e294f737f4c.vhd when simulating
-- the core, cntr_11_0_86806e294f737f4c. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_86806e294f737f4c IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_86806e294f737f4c;

ARCHITECTURE cntr_11_0_86806e294f737f4c_a OF cntr_11_0_86806e294f737f4c IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_86806e294f737f4c
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_86806e294f737f4c USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_86806e294f737f4c
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_86806e294f737f4c_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_bcc28bfecf25caff.vhd when simulating
-- the core, cntr_11_0_bcc28bfecf25caff. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_bcc28bfecf25caff IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END cntr_11_0_bcc28bfecf25caff;

ARCHITECTURE cntr_11_0_bcc28bfecf25caff_a OF cntr_11_0_bcc28bfecf25caff IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_bcc28bfecf25caff
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_bcc28bfecf25caff USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 3,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_bcc28bfecf25caff
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_bcc28bfecf25caff_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_d24951bef2f0cdc9.vhd when simulating
-- the core, cntr_11_0_d24951bef2f0cdc9. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_d24951bef2f0cdc9 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END cntr_11_0_d24951bef2f0cdc9;

ARCHITECTURE cntr_11_0_d24951bef2f0cdc9_a OF cntr_11_0_d24951bef2f0cdc9 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_d24951bef2f0cdc9
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_d24951bef2f0cdc9 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 7,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_d24951bef2f0cdc9
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_d24951bef2f0cdc9_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_d66925a45384983e.vhd when simulating
-- the core, cntr_11_0_d66925a45384983e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_d66925a45384983e IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END cntr_11_0_d66925a45384983e;

ARCHITECTURE cntr_11_0_d66925a45384983e_a OF cntr_11_0_d66925a45384983e IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_d66925a45384983e
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_d66925a45384983e USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "1",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 9,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_d66925a45384983e
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_d66925a45384983e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_f068fb73312ae1e5.vhd when simulating
-- the core, cntr_11_0_f068fb73312ae1e5. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_f068fb73312ae1e5 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END cntr_11_0_f068fb73312ae1e5;

ARCHITECTURE cntr_11_0_f068fb73312ae1e5_a OF cntr_11_0_f068fb73312ae1e5 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_f068fb73312ae1e5
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_f068fb73312ae1e5 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 6,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_f068fb73312ae1e5
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_f068fb73312ae1e5_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_134e91999cae8947.vhd when simulating
-- the core, dmg_72_134e91999cae8947. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_134e91999cae8947 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END dmg_72_134e91999cae8947;

ARCHITECTURE dmg_72_134e91999cae8947_a OF dmg_72_134e91999cae8947 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_134e91999cae8947
  PORT (
    a : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_134e91999cae8947 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 8,
      c_default_data => "0",
      c_depth => 256,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_134e91999cae8947.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 32
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_134e91999cae8947
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_134e91999cae8947_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_140171b6b191950b.vhd when simulating
-- the core, dmg_72_140171b6b191950b. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_140171b6b191950b IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_140171b6b191950b;

ARCHITECTURE dmg_72_140171b6b191950b_a OF dmg_72_140171b6b191950b IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_140171b6b191950b
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_140171b6b191950b USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 9,
      c_default_data => "0",
      c_depth => 512,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_140171b6b191950b.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_140171b6b191950b
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_140171b6b191950b_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_28ec6cac12d9767d.vhd when simulating
-- the core, dmg_72_28ec6cac12d9767d. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_28ec6cac12d9767d IS
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END dmg_72_28ec6cac12d9767d;

ARCHITECTURE dmg_72_28ec6cac12d9767d_a OF dmg_72_28ec6cac12d9767d IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_28ec6cac12d9767d
  PORT (
    a : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
    clk : IN STD_LOGIC;
    qspo_ce : IN STD_LOGIC;
    qspo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_28ec6cac12d9767d USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 9,
      c_default_data => "0",
      c_depth => 512,
      c_family => "virtex6",
      c_has_clk => 1,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 1,
      c_has_qspo_ce => 1,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 0,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_28ec6cac12d9767d.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 16
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_28ec6cac12d9767d
  PORT MAP (
    a => a,
    clk => clk,
    qspo_ce => qspo_ce,
    qspo => qspo
  );
-- synthesis translate_on

END dmg_72_28ec6cac12d9767d_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file dmg_72_5efcdb43c0011b51.vhd when simulating
-- the core, dmg_72_5efcdb43c0011b51. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY dmg_72_5efcdb43c0011b51 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END dmg_72_5efcdb43c0011b51;

ARCHITECTURE dmg_72_5efcdb43c0011b51_a OF dmg_72_5efcdb43c0011b51 IS
-- synthesis translate_off
COMPONENT wrapped_dmg_72_5efcdb43c0011b51
  PORT (
    a : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    spo : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_dmg_72_5efcdb43c0011b51 USE ENTITY XilinxCoreLib.dist_mem_gen_v7_2(behavioral)
    GENERIC MAP (
      c_addr_width => 6,
      c_default_data => "0",
      c_depth => 64,
      c_family => "virtex6",
      c_has_clk => 0,
      c_has_d => 0,
      c_has_dpo => 0,
      c_has_dpra => 0,
      c_has_i_ce => 0,
      c_has_qdpo => 0,
      c_has_qdpo_ce => 0,
      c_has_qdpo_clk => 0,
      c_has_qdpo_rst => 0,
      c_has_qdpo_srst => 0,
      c_has_qspo => 0,
      c_has_qspo_ce => 0,
      c_has_qspo_rst => 0,
      c_has_qspo_srst => 0,
      c_has_spo => 1,
      c_has_spra => 0,
      c_has_we => 0,
      c_mem_init_file => "dmg_72_5efcdb43c0011b51.mif",
      c_mem_type => 0,
      c_parser_type => 1,
      c_pipeline_stages => 0,
      c_qce_joined => 0,
      c_qualify_we => 0,
      c_read_mif => 1,
      c_reg_a_d_inputs => 0,
      c_reg_dpra_input => 0,
      c_sync_enable => 1,
      c_width => 7
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_dmg_72_5efcdb43c0011b51
  PORT MAP (
    a => a,
    spo => spo
  );
-- synthesis translate_on

END dmg_72_5efcdb43c0011b51_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file fifo_fg92_6a1156e8dc43a711.vhd when simulating
-- the core, fifo_fg92_6a1156e8dc43a711. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY fifo_fg92_6a1156e8dc43a711 IS
  PORT (
    clk : IN STD_LOGIC;
    srst : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC;
    data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END fifo_fg92_6a1156e8dc43a711;

ARCHITECTURE fifo_fg92_6a1156e8dc43a711_a OF fifo_fg92_6a1156e8dc43a711 IS
-- synthesis translate_off
COMPONENT wrapped_fifo_fg92_6a1156e8dc43a711
  PORT (
    clk : IN STD_LOGIC;
    srst : IN STD_LOGIC;
    din : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    wr_en : IN STD_LOGIC;
    rd_en : IN STD_LOGIC;
    dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    full : OUT STD_LOGIC;
    empty : OUT STD_LOGIC;
    data_count : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_fifo_fg92_6a1156e8dc43a711 USE ENTITY XilinxCoreLib.fifo_generator_v9_3(behavioral)
    GENERIC MAP (
      c_add_ngc_constraint => 0,
      c_application_type_axis => 0,
      c_application_type_rach => 0,
      c_application_type_rdch => 0,
      c_application_type_wach => 0,
      c_application_type_wdch => 0,
      c_application_type_wrch => 0,
      c_axi_addr_width => 32,
      c_axi_aruser_width => 1,
      c_axi_awuser_width => 1,
      c_axi_buser_width => 1,
      c_axi_data_width => 64,
      c_axi_id_width => 4,
      c_axi_ruser_width => 1,
      c_axi_type => 0,
      c_axi_wuser_width => 1,
      c_axis_tdata_width => 64,
      c_axis_tdest_width => 4,
      c_axis_tid_width => 8,
      c_axis_tkeep_width => 4,
      c_axis_tstrb_width => 4,
      c_axis_tuser_width => 4,
      c_axis_type => 0,
      c_common_clock => 1,
      c_count_type => 0,
      c_data_count_width => 8,
      c_default_value => "BlankString",
      c_din_width => 32,
      c_din_width_axis => 1,
      c_din_width_rach => 32,
      c_din_width_rdch => 64,
      c_din_width_wach => 32,
      c_din_width_wdch => 64,
      c_din_width_wrch => 2,
      c_dout_rst_val => "0",
      c_dout_width => 32,
      c_enable_rlocs => 0,
      c_enable_rst_sync => 1,
      c_error_injection_type => 0,
      c_error_injection_type_axis => 0,
      c_error_injection_type_rach => 0,
      c_error_injection_type_rdch => 0,
      c_error_injection_type_wach => 0,
      c_error_injection_type_wdch => 0,
      c_error_injection_type_wrch => 0,
      c_family => "virtex6",
      c_full_flags_rst_val => 0,
      c_has_almost_empty => 0,
      c_has_almost_full => 0,
      c_has_axi_aruser => 0,
      c_has_axi_awuser => 0,
      c_has_axi_buser => 0,
      c_has_axi_rd_channel => 0,
      c_has_axi_ruser => 0,
      c_has_axi_wr_channel => 0,
      c_has_axi_wuser => 0,
      c_has_axis_tdata => 0,
      c_has_axis_tdest => 0,
      c_has_axis_tid => 0,
      c_has_axis_tkeep => 0,
      c_has_axis_tlast => 0,
      c_has_axis_tready => 1,
      c_has_axis_tstrb => 0,
      c_has_axis_tuser => 0,
      c_has_backup => 0,
      c_has_data_count => 1,
      c_has_data_counts_axis => 0,
      c_has_data_counts_rach => 0,
      c_has_data_counts_rdch => 0,
      c_has_data_counts_wach => 0,
      c_has_data_counts_wdch => 0,
      c_has_data_counts_wrch => 0,
      c_has_int_clk => 0,
      c_has_master_ce => 0,
      c_has_meminit_file => 0,
      c_has_overflow => 0,
      c_has_prog_flags_axis => 0,
      c_has_prog_flags_rach => 0,
      c_has_prog_flags_rdch => 0,
      c_has_prog_flags_wach => 0,
      c_has_prog_flags_wdch => 0,
      c_has_prog_flags_wrch => 0,
      c_has_rd_data_count => 0,
      c_has_rd_rst => 0,
      c_has_rst => 0,
      c_has_slave_ce => 0,
      c_has_srst => 1,
      c_has_underflow => 0,
      c_has_valid => 0,
      c_has_wr_ack => 0,
      c_has_wr_data_count => 0,
      c_has_wr_rst => 0,
      c_implementation_type => 0,
      c_implementation_type_axis => 1,
      c_implementation_type_rach => 1,
      c_implementation_type_rdch => 1,
      c_implementation_type_wach => 1,
      c_implementation_type_wdch => 1,
      c_implementation_type_wrch => 1,
      c_init_wr_pntr_val => 0,
      c_interface_type => 0,
      c_memory_type => 1,
      c_mif_file_name => "BlankString",
      c_msgon_val => 1,
      c_optimization_mode => 0,
      c_overflow_low => 0,
      c_preload_latency => 2,
      c_preload_regs => 1,
      c_prim_fifo_type => "512x36",
      c_prog_empty_thresh_assert_val => 2,
      c_prog_empty_thresh_assert_val_axis => 1022,
      c_prog_empty_thresh_assert_val_rach => 1022,
      c_prog_empty_thresh_assert_val_rdch => 1022,
      c_prog_empty_thresh_assert_val_wach => 1022,
      c_prog_empty_thresh_assert_val_wdch => 1022,
      c_prog_empty_thresh_assert_val_wrch => 1022,
      c_prog_empty_thresh_negate_val => 3,
      c_prog_empty_type => 0,
      c_prog_empty_type_axis => 0,
      c_prog_empty_type_rach => 0,
      c_prog_empty_type_rdch => 0,
      c_prog_empty_type_wach => 0,
      c_prog_empty_type_wdch => 0,
      c_prog_empty_type_wrch => 0,
      c_prog_full_thresh_assert_val => 254,
      c_prog_full_thresh_assert_val_axis => 1023,
      c_prog_full_thresh_assert_val_rach => 1023,
      c_prog_full_thresh_assert_val_rdch => 1023,
      c_prog_full_thresh_assert_val_wach => 1023,
      c_prog_full_thresh_assert_val_wdch => 1023,
      c_prog_full_thresh_assert_val_wrch => 1023,
      c_prog_full_thresh_negate_val => 253,
      c_prog_full_type => 0,
      c_prog_full_type_axis => 0,
      c_prog_full_type_rach => 0,
      c_prog_full_type_rdch => 0,
      c_prog_full_type_wach => 0,
      c_prog_full_type_wdch => 0,
      c_prog_full_type_wrch => 0,
      c_rach_type => 0,
      c_rd_data_count_width => 8,
      c_rd_depth => 256,
      c_rd_freq => 1,
      c_rd_pntr_width => 8,
      c_rdch_type => 0,
      c_reg_slice_mode_axis => 0,
      c_reg_slice_mode_rach => 0,
      c_reg_slice_mode_rdch => 0,
      c_reg_slice_mode_wach => 0,
      c_reg_slice_mode_wdch => 0,
      c_reg_slice_mode_wrch => 0,
      c_synchronizer_stage => 2,
      c_underflow_low => 0,
      c_use_common_overflow => 0,
      c_use_common_underflow => 0,
      c_use_default_settings => 0,
      c_use_dout_rst => 1,
      c_use_ecc => 0,
      c_use_ecc_axis => 0,
      c_use_ecc_rach => 0,
      c_use_ecc_rdch => 0,
      c_use_ecc_wach => 0,
      c_use_ecc_wdch => 0,
      c_use_ecc_wrch => 0,
      c_use_embedded_reg => 1,
      c_use_fifo16_flags => 0,
      c_use_fwft_data_count => 0,
      c_valid_low => 0,
      c_wach_type => 0,
      c_wdch_type => 0,
      c_wr_ack_low => 0,
      c_wr_data_count_width => 8,
      c_wr_depth => 256,
      c_wr_depth_axis => 1024,
      c_wr_depth_rach => 16,
      c_wr_depth_rdch => 1024,
      c_wr_depth_wach => 16,
      c_wr_depth_wdch => 1024,
      c_wr_depth_wrch => 16,
      c_wr_freq => 1,
      c_wr_pntr_width => 8,
      c_wr_pntr_width_axis => 10,
      c_wr_pntr_width_rach => 4,
      c_wr_pntr_width_rdch => 10,
      c_wr_pntr_width_wach => 4,
      c_wr_pntr_width_wdch => 10,
      c_wr_pntr_width_wrch => 4,
      c_wr_response_latency => 1,
      c_wrch_type => 0
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_fifo_fg92_6a1156e8dc43a711
  PORT MAP (
    clk => clk,
    srst => srst,
    din => din,
    wr_en => wr_en,
    rd_en => rd_en,
    dout => dout,
    full => full,
    empty => empty,
    data_count => data_count
  );
-- synthesis translate_on

END fifo_fg92_6a1156e8dc43a711_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_414c0fa5acc33f35.vhd when simulating
-- the core, mult_11_2_414c0fa5acc33f35. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_414c0fa5acc33f35 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END mult_11_2_414c0fa5acc33f35;

ARCHITECTURE mult_11_2_414c0fa5acc33f35_a OF mult_11_2_414c0fa5acc33f35 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_414c0fa5acc33f35
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_414c0fa5acc33f35 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 0,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_zero_detect => 0,
      c_latency => 0,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 31,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_414c0fa5acc33f35
  PORT MAP (
    a => a,
    b => b,
    p => p
  );
-- synthesis translate_on

END mult_11_2_414c0fa5acc33f35_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2013 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_f2bb5a57782af7d9.vhd when simulating
-- the core, mult_11_2_f2bb5a57782af7d9. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_f2bb5a57782af7d9 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END mult_11_2_f2bb5a57782af7d9;

ARCHITECTURE mult_11_2_f2bb5a57782af7d9_a OF mult_11_2_f2bb5a57782af7d9 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_f2bb5a57782af7d9
  PORT (
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_f2bb5a57782af7d9 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 0,
      c_a_width => 16,
      c_b_type => 1,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_zero_detect => 0,
      c_latency => 0,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 31,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_f2bb5a57782af7d9
  PORT MAP (
    a => a,
    b => b,
    p => p
  );
-- synthesis translate_on

END mult_11_2_f2bb5a57782af7d9_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2012 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: P.49d
--  \   \         Application: netgen
--  /   /         Filename: xfft_v8_0_6e4d6522fcd78ca0.vhd
-- /___/   /\     Timestamp: Mon Jul 29 22:38:54 2013
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -w -sim -ofmt vhdl S:/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c48e2efa8eb3b3387/tmp/_cg/xfft_v8_0_6e4d6522fcd78ca0.ngc S:/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c48e2efa8eb3b3387/tmp/_cg/xfft_v8_0_6e4d6522fcd78ca0.vhd 
-- Device	: 6vlx240tff1156-2
-- Input file	: S:/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c48e2efa8eb3b3387/tmp/_cg/xfft_v8_0_6e4d6522fcd78ca0.ngc
-- Output file	: S:/murphpo/AppData/Local/Temp/sysgentmp-murphpo/cg_wk/c48e2efa8eb3b3387/tmp/_cg/xfft_v8_0_6e4d6522fcd78ca0.vhd
-- # of Entities	: 1
-- Design Name	: xfft_v8_0_6e4d6522fcd78ca0
-- Xilinx	: s:\xilinx\14.4\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity xfft_v8_0_6e4d6522fcd78ca0 is
  port (
    aclk : in STD_LOGIC := 'X'; 
    aclken : in STD_LOGIC := 'X'; 
    aresetn : in STD_LOGIC := 'X'; 
    s_axis_config_tvalid : in STD_LOGIC := 'X'; 
    s_axis_data_tvalid : in STD_LOGIC := 'X'; 
    s_axis_data_tlast : in STD_LOGIC := 'X'; 
    m_axis_data_tready : in STD_LOGIC := 'X'; 
    m_axis_status_tready : in STD_LOGIC := 'X'; 
    s_axis_config_tready : out STD_LOGIC; 
    s_axis_data_tready : out STD_LOGIC; 
    m_axis_data_tvalid : out STD_LOGIC; 
    m_axis_data_tlast : out STD_LOGIC; 
    m_axis_status_tvalid : out STD_LOGIC; 
    event_frame_started : out STD_LOGIC; 
    event_tlast_unexpected : out STD_LOGIC; 
    event_tlast_missing : out STD_LOGIC; 
    event_fft_overflow : out STD_LOGIC; 
    event_status_channel_halt : out STD_LOGIC; 
    event_data_in_channel_halt : out STD_LOGIC; 
    event_data_out_channel_halt : out STD_LOGIC; 
    s_axis_config_tdata : in STD_LOGIC_VECTOR ( 15 downto 0 ); 
    s_axis_data_tdata : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    m_axis_data_tdata : out STD_LOGIC_VECTOR ( 31 downto 0 ); 
    m_axis_data_tuser : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    m_axis_status_tdata : out STD_LOGIC_VECTOR ( 7 downto 0 ) 
  );
end xfft_v8_0_6e4d6522fcd78ca0;

architecture STRUCTURE of xfft_v8_0_6e4d6522fcd78ca0 is
  signal NlwRenamedSig_OI_m_axis_data_tuser_10_Q : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_data_tuser_8_Q : STD_LOGIC; 
  signal NlwRenamedSig_OI_s_axis_config_tready : STD_LOGIC; 
  signal NlwRenamedSig_OI_s_axis_data_tready : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_data_tvalid : STD_LOGIC; 
  signal NlwRenamedSig_OI_m_axis_status_tvalid : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_frame_started : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_tlast_missing : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_fft_overflow : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_status_channel_halt : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_data_in_channel_halt : STD_LOGIC; 
  signal NlwRenamedSig_OI_event_data_out_channel_halt : STD_LOGIC; 
  signal blk00000001_sig000001be : STD_LOGIC; 
  signal blk00000001_sig000001bd : STD_LOGIC; 
  signal blk00000001_sig000001bc : STD_LOGIC; 
  signal blk00000001_sig000001bb : STD_LOGIC; 
  signal blk00000001_sig000001ba : STD_LOGIC; 
  signal blk00000001_sig000001b9 : STD_LOGIC; 
  signal blk00000001_sig000001b8 : STD_LOGIC; 
  signal blk00000001_sig000001b7 : STD_LOGIC; 
  signal blk00000001_sig000001b6 : STD_LOGIC; 
  signal blk00000001_sig000001b5 : STD_LOGIC; 
  signal blk00000001_sig000001b4 : STD_LOGIC; 
  signal blk00000001_sig000001b3 : STD_LOGIC; 
  signal blk00000001_sig000001b2 : STD_LOGIC; 
  signal blk00000001_sig000001b1 : STD_LOGIC; 
  signal blk00000001_sig000001b0 : STD_LOGIC; 
  signal blk00000001_sig000001af : STD_LOGIC; 
  signal blk00000001_sig000001ae : STD_LOGIC; 
  signal blk00000001_sig000001ad : STD_LOGIC; 
  signal blk00000001_sig000001ac : STD_LOGIC; 
  signal blk00000001_sig000001ab : STD_LOGIC; 
  signal blk00000001_sig000001aa : STD_LOGIC; 
  signal blk00000001_sig000001a9 : STD_LOGIC; 
  signal blk00000001_sig000001a8 : STD_LOGIC; 
  signal blk00000001_sig000001a7 : STD_LOGIC; 
  signal blk00000001_sig000001a6 : STD_LOGIC; 
  signal blk00000001_sig000001a5 : STD_LOGIC; 
  signal blk00000001_sig000001a4 : STD_LOGIC; 
  signal blk00000001_sig000001a3 : STD_LOGIC; 
  signal blk00000001_sig000001a2 : STD_LOGIC; 
  signal blk00000001_sig000001a1 : STD_LOGIC; 
  signal blk00000001_sig000001a0 : STD_LOGIC; 
  signal blk00000001_sig0000019f : STD_LOGIC; 
  signal blk00000001_sig0000019e : STD_LOGIC; 
  signal blk00000001_sig0000019d : STD_LOGIC; 
  signal blk00000001_sig0000019c : STD_LOGIC; 
  signal blk00000001_sig0000019b : STD_LOGIC; 
  signal blk00000001_sig0000019a : STD_LOGIC; 
  signal blk00000001_sig00000199 : STD_LOGIC; 
  signal blk00000001_sig00000198 : STD_LOGIC; 
  signal blk00000001_sig00000197 : STD_LOGIC; 
  signal blk00000001_sig00000196 : STD_LOGIC; 
  signal blk00000001_sig00000195 : STD_LOGIC; 
  signal blk00000001_sig00000194 : STD_LOGIC; 
  signal blk00000001_sig00000193 : STD_LOGIC; 
  signal blk00000001_sig00000192 : STD_LOGIC; 
  signal blk00000001_sig00000191 : STD_LOGIC; 
  signal blk00000001_sig00000190 : STD_LOGIC; 
  signal blk00000001_sig0000018f : STD_LOGIC; 
  signal blk00000001_sig0000018e : STD_LOGIC; 
  signal blk00000001_sig0000018d : STD_LOGIC; 
  signal blk00000001_sig0000018c : STD_LOGIC; 
  signal blk00000001_sig0000018b : STD_LOGIC; 
  signal blk00000001_sig0000018a : STD_LOGIC; 
  signal blk00000001_sig00000189 : STD_LOGIC; 
  signal blk00000001_sig00000188 : STD_LOGIC; 
  signal blk00000001_sig00000187 : STD_LOGIC; 
  signal blk00000001_sig00000186 : STD_LOGIC; 
  signal blk00000001_sig00000185 : STD_LOGIC; 
  signal blk00000001_sig00000184 : STD_LOGIC; 
  signal blk00000001_sig00000183 : STD_LOGIC; 
  signal blk00000001_sig00000182 : STD_LOGIC; 
  signal blk00000001_sig00000181 : STD_LOGIC; 
  signal blk00000001_sig00000180 : STD_LOGIC; 
  signal blk00000001_sig0000017f : STD_LOGIC; 
  signal blk00000001_sig0000017e : STD_LOGIC; 
  signal blk00000001_sig0000017d : STD_LOGIC; 
  signal blk00000001_sig0000017c : STD_LOGIC; 
  signal blk00000001_sig0000017b : STD_LOGIC; 
  signal blk00000001_sig0000017a : STD_LOGIC; 
  signal blk00000001_sig00000179 : STD_LOGIC; 
  signal blk00000001_sig00000178 : STD_LOGIC; 
  signal blk00000001_sig00000177 : STD_LOGIC; 
  signal blk00000001_sig00000176 : STD_LOGIC; 
  signal blk00000001_sig00000175 : STD_LOGIC; 
  signal blk00000001_sig00000174 : STD_LOGIC; 
  signal blk00000001_sig00000173 : STD_LOGIC; 
  signal blk00000001_sig00000172 : STD_LOGIC; 
  signal blk00000001_sig00000171 : STD_LOGIC; 
  signal blk00000001_sig00000170 : STD_LOGIC; 
  signal blk00000001_sig0000016f : STD_LOGIC; 
  signal blk00000001_sig0000016e : STD_LOGIC; 
  signal blk00000001_sig0000016d : STD_LOGIC; 
  signal blk00000001_sig0000016c : STD_LOGIC; 
  signal blk00000001_sig0000016b : STD_LOGIC; 
  signal blk00000001_sig0000016a : STD_LOGIC; 
  signal blk00000001_sig00000169 : STD_LOGIC; 
  signal blk00000001_sig00000168 : STD_LOGIC; 
  signal blk00000001_sig00000167 : STD_LOGIC; 
  signal blk00000001_sig00000166 : STD_LOGIC; 
  signal blk00000001_sig00000165 : STD_LOGIC; 
  signal blk00000001_sig00000164 : STD_LOGIC; 
  signal blk00000001_sig00000163 : STD_LOGIC; 
  signal blk00000001_sig00000162 : STD_LOGIC; 
  signal blk00000001_sig00000161 : STD_LOGIC; 
  signal blk00000001_sig00000160 : STD_LOGIC; 
  signal blk00000001_sig0000015f : STD_LOGIC; 
  signal blk00000001_sig0000015e : STD_LOGIC; 
  signal blk00000001_sig0000015d : STD_LOGIC; 
  signal blk00000001_sig0000015c : STD_LOGIC; 
  signal blk00000001_sig0000015b : STD_LOGIC; 
  signal blk00000001_sig0000015a : STD_LOGIC; 
  signal blk00000001_sig00000159 : STD_LOGIC; 
  signal blk00000001_sig00000158 : STD_LOGIC; 
  signal blk00000001_sig00000157 : STD_LOGIC; 
  signal blk00000001_sig00000156 : STD_LOGIC; 
  signal blk00000001_sig00000155 : STD_LOGIC; 
  signal blk00000001_sig00000154 : STD_LOGIC; 
  signal blk00000001_sig00000153 : STD_LOGIC; 
  signal blk00000001_sig00000152 : STD_LOGIC; 
  signal blk00000001_sig00000151 : STD_LOGIC; 
  signal blk00000001_sig00000150 : STD_LOGIC; 
  signal blk00000001_sig0000014f : STD_LOGIC; 
  signal blk00000001_sig0000014e : STD_LOGIC; 
  signal blk00000001_sig0000014d : STD_LOGIC; 
  signal blk00000001_sig0000014c : STD_LOGIC; 
  signal blk00000001_sig0000014b : STD_LOGIC; 
  signal blk00000001_sig0000014a : STD_LOGIC; 
  signal blk00000001_sig00000149 : STD_LOGIC; 
  signal blk00000001_sig00000148 : STD_LOGIC; 
  signal blk00000001_sig00000147 : STD_LOGIC; 
  signal blk00000001_sig00000146 : STD_LOGIC; 
  signal blk00000001_sig00000145 : STD_LOGIC; 
  signal blk00000001_sig00000144 : STD_LOGIC; 
  signal blk00000001_sig00000143 : STD_LOGIC; 
  signal blk00000001_sig00000142 : STD_LOGIC; 
  signal blk00000001_sig00000141 : STD_LOGIC; 
  signal blk00000001_sig00000140 : STD_LOGIC; 
  signal blk00000001_sig0000013f : STD_LOGIC; 
  signal blk00000001_sig0000013e : STD_LOGIC; 
  signal blk00000001_sig0000013d : STD_LOGIC; 
  signal blk00000001_sig0000013c : STD_LOGIC; 
  signal blk00000001_sig0000013b : STD_LOGIC; 
  signal blk00000001_sig0000013a : STD_LOGIC; 
  signal blk00000001_sig00000139 : STD_LOGIC; 
  signal blk00000001_sig00000138 : STD_LOGIC; 
  signal blk00000001_sig00000137 : STD_LOGIC; 
  signal blk00000001_sig00000136 : STD_LOGIC; 
  signal blk00000001_sig00000135 : STD_LOGIC; 
  signal blk00000001_sig00000134 : STD_LOGIC; 
  signal blk00000001_sig00000133 : STD_LOGIC; 
  signal blk00000001_sig00000132 : STD_LOGIC; 
  signal blk00000001_sig00000131 : STD_LOGIC; 
  signal blk00000001_sig00000130 : STD_LOGIC; 
  signal blk00000001_sig0000012f : STD_LOGIC; 
  signal blk00000001_sig0000012e : STD_LOGIC; 
  signal blk00000001_sig0000012d : STD_LOGIC; 
  signal blk00000001_sig0000012c : STD_LOGIC; 
  signal blk00000001_sig0000012b : STD_LOGIC; 
  signal blk00000001_sig0000012a : STD_LOGIC; 
  signal blk00000001_sig00000129 : STD_LOGIC; 
  signal blk00000001_sig00000128 : STD_LOGIC; 
  signal blk00000001_sig00000127 : STD_LOGIC; 
  signal blk00000001_sig00000126 : STD_LOGIC; 
  signal blk00000001_sig00000125 : STD_LOGIC; 
  signal blk00000001_sig00000124 : STD_LOGIC; 
  signal blk00000001_sig00000123 : STD_LOGIC; 
  signal blk00000001_sig00000122 : STD_LOGIC; 
  signal blk00000001_sig00000121 : STD_LOGIC; 
  signal blk00000001_sig00000120 : STD_LOGIC; 
  signal blk00000001_sig0000011f : STD_LOGIC; 
  signal blk00000001_sig0000011e : STD_LOGIC; 
  signal blk00000001_sig0000011d : STD_LOGIC; 
  signal blk00000001_sig0000011c : STD_LOGIC; 
  signal blk00000001_sig0000011b : STD_LOGIC; 
  signal blk00000001_sig0000011a : STD_LOGIC; 
  signal blk00000001_sig00000119 : STD_LOGIC; 
  signal blk00000001_sig00000118 : STD_LOGIC; 
  signal blk00000001_sig00000117 : STD_LOGIC; 
  signal blk00000001_sig00000116 : STD_LOGIC; 
  signal blk00000001_sig00000115 : STD_LOGIC; 
  signal blk00000001_sig00000114 : STD_LOGIC; 
  signal blk00000001_sig00000113 : STD_LOGIC; 
  signal blk00000001_sig00000112 : STD_LOGIC; 
  signal blk00000001_sig00000111 : STD_LOGIC; 
  signal blk00000001_sig00000110 : STD_LOGIC; 
  signal blk00000001_sig0000010f : STD_LOGIC; 
  signal blk00000001_sig0000010e : STD_LOGIC; 
  signal blk00000001_sig0000010d : STD_LOGIC; 
  signal blk00000001_sig0000010c : STD_LOGIC; 
  signal blk00000001_sig0000010b : STD_LOGIC; 
  signal blk00000001_sig0000010a : STD_LOGIC; 
  signal blk00000001_sig00000109 : STD_LOGIC; 
  signal blk00000001_sig00000108 : STD_LOGIC; 
  signal blk00000001_sig00000107 : STD_LOGIC; 
  signal blk00000001_sig00000106 : STD_LOGIC; 
  signal blk00000001_sig00000105 : STD_LOGIC; 
  signal blk00000001_sig00000104 : STD_LOGIC; 
  signal blk00000001_sig00000103 : STD_LOGIC; 
  signal blk00000001_sig00000102 : STD_LOGIC; 
  signal blk00000001_sig00000101 : STD_LOGIC; 
  signal blk00000001_sig00000100 : STD_LOGIC; 
  signal blk00000001_sig000000ff : STD_LOGIC; 
  signal blk00000001_sig000000fe : STD_LOGIC; 
  signal blk00000001_sig000000fd : STD_LOGIC; 
  signal blk00000001_sig000000fc : STD_LOGIC; 
  signal blk00000001_sig000000fb : STD_LOGIC; 
  signal blk00000001_sig000000fa : STD_LOGIC; 
  signal blk00000001_sig000000f9 : STD_LOGIC; 
  signal blk00000001_sig000000f8 : STD_LOGIC; 
  signal blk00000001_sig000000f7 : STD_LOGIC; 
  signal blk00000001_sig000000f6 : STD_LOGIC; 
  signal blk00000001_sig000000f5 : STD_LOGIC; 
  signal blk00000001_sig000000f4 : STD_LOGIC; 
  signal blk00000001_sig000000f3 : STD_LOGIC; 
  signal blk00000001_sig000000f2 : STD_LOGIC; 
  signal blk00000001_sig000000f1 : STD_LOGIC; 
  signal blk00000001_sig000000f0 : STD_LOGIC; 
  signal blk00000001_sig000000ef : STD_LOGIC; 
  signal blk00000001_sig000000ee : STD_LOGIC; 
  signal blk00000001_sig000000ed : STD_LOGIC; 
  signal blk00000001_sig000000ec : STD_LOGIC; 
  signal blk00000001_sig000000eb : STD_LOGIC; 
  signal blk00000001_sig000000ea : STD_LOGIC; 
  signal blk00000001_sig000000e9 : STD_LOGIC; 
  signal blk00000001_sig000000e8 : STD_LOGIC; 
  signal blk00000001_sig000000e7 : STD_LOGIC; 
  signal blk00000001_sig000000e6 : STD_LOGIC; 
  signal blk00000001_sig000000e5 : STD_LOGIC; 
  signal blk00000001_sig000000e4 : STD_LOGIC; 
  signal blk00000001_sig000000e3 : STD_LOGIC; 
  signal blk00000001_sig000000e2 : STD_LOGIC; 
  signal blk00000001_sig000000e1 : STD_LOGIC; 
  signal blk00000001_sig000000e0 : STD_LOGIC; 
  signal blk00000001_sig000000df : STD_LOGIC; 
  signal blk00000001_sig000000de : STD_LOGIC; 
  signal blk00000001_sig000000dd : STD_LOGIC; 
  signal blk00000001_sig000000dc : STD_LOGIC; 
  signal blk00000001_sig000000db : STD_LOGIC; 
  signal blk00000001_sig000000da : STD_LOGIC; 
  signal blk00000001_sig000000d9 : STD_LOGIC; 
  signal blk00000001_sig000000d8 : STD_LOGIC; 
  signal blk00000001_sig000000d7 : STD_LOGIC; 
  signal blk00000001_sig000000d6 : STD_LOGIC; 
  signal blk00000001_sig000000d5 : STD_LOGIC; 
  signal blk00000001_sig000000d4 : STD_LOGIC; 
  signal blk00000001_sig000000d3 : STD_LOGIC; 
  signal blk00000001_sig000000d2 : STD_LOGIC; 
  signal blk00000001_sig000000d1 : STD_LOGIC; 
  signal blk00000001_sig000000d0 : STD_LOGIC; 
  signal blk00000001_sig000000cf : STD_LOGIC; 
  signal blk00000001_sig000000ce : STD_LOGIC; 
  signal blk00000001_sig000000cd : STD_LOGIC; 
  signal blk00000001_sig000000cb : STD_LOGIC; 
  signal blk00000001_sig000000ca : STD_LOGIC; 
  signal blk00000001_sig000000c9 : STD_LOGIC; 
  signal blk00000001_sig000000c8 : STD_LOGIC; 
  signal blk00000001_sig000000c7 : STD_LOGIC; 
  signal blk00000001_sig000000c6 : STD_LOGIC; 
  signal blk00000001_sig000000c5 : STD_LOGIC; 
  signal blk00000001_sig000000c4 : STD_LOGIC; 
  signal blk00000001_sig000000c3 : STD_LOGIC; 
  signal blk00000001_sig000000c2 : STD_LOGIC; 
  signal blk00000001_sig000000c1 : STD_LOGIC; 
  signal blk00000001_sig000000c0 : STD_LOGIC; 
  signal blk00000001_sig000000bf : STD_LOGIC; 
  signal blk00000001_sig000000be : STD_LOGIC; 
  signal blk00000001_sig000000bd : STD_LOGIC; 
  signal blk00000001_sig000000bc : STD_LOGIC; 
  signal blk00000001_sig000000bb : STD_LOGIC; 
  signal blk00000001_sig000000ba : STD_LOGIC; 
  signal blk00000001_sig000000b9 : STD_LOGIC; 
  signal blk00000001_sig000000b8 : STD_LOGIC; 
  signal blk00000001_sig000000b7 : STD_LOGIC; 
  signal blk00000001_sig000000b6 : STD_LOGIC; 
  signal blk00000001_sig000000b5 : STD_LOGIC; 
  signal blk00000001_sig000000b4 : STD_LOGIC; 
  signal blk00000001_sig000000b3 : STD_LOGIC; 
  signal blk00000001_sig000000b2 : STD_LOGIC; 
  signal blk00000001_sig000000b1 : STD_LOGIC; 
  signal blk00000001_sig000000b0 : STD_LOGIC; 
  signal blk00000001_sig000000af : STD_LOGIC; 
  signal blk00000001_sig000000ae : STD_LOGIC; 
  signal blk00000001_sig000000ad : STD_LOGIC; 
  signal blk00000001_sig000000ac : STD_LOGIC; 
  signal blk00000001_sig000000ab : STD_LOGIC; 
  signal blk00000001_sig000000aa : STD_LOGIC; 
  signal blk00000001_sig000000a9 : STD_LOGIC; 
  signal blk00000001_sig000000a8 : STD_LOGIC; 
  signal blk00000001_sig000000a7 : STD_LOGIC; 
  signal blk00000001_sig000000a6 : STD_LOGIC; 
  signal blk00000001_sig000000a5 : STD_LOGIC; 
  signal blk00000001_sig000000a4 : STD_LOGIC; 
  signal blk00000001_sig000000a3 : STD_LOGIC; 
  signal blk00000001_sig000000a2 : STD_LOGIC; 
  signal blk00000001_sig000000a1 : STD_LOGIC; 
  signal blk00000001_sig000000a0 : STD_LOGIC; 
  signal blk00000001_sig0000009f : STD_LOGIC; 
  signal blk00000001_sig0000009e : STD_LOGIC; 
  signal blk00000001_sig0000009d : STD_LOGIC; 
  signal blk00000001_sig0000009c : STD_LOGIC; 
  signal blk00000001_sig0000009b : STD_LOGIC; 
  signal blk00000001_sig0000009a : STD_LOGIC; 
  signal blk00000001_sig00000099 : STD_LOGIC; 
  signal blk00000001_sig00000098 : STD_LOGIC; 
  signal blk00000001_sig00000097 : STD_LOGIC; 
  signal blk00000001_sig00000096 : STD_LOGIC; 
  signal blk00000001_sig00000089 : STD_LOGIC; 
  signal blk00000001_sig00000088 : STD_LOGIC; 
  signal blk00000001_sig00000087 : STD_LOGIC; 
  signal blk00000001_sig00000086 : STD_LOGIC; 
  signal blk00000001_sig00000085 : STD_LOGIC; 
  signal blk00000001_sig00000084 : STD_LOGIC; 
  signal blk00000001_sig00000083 : STD_LOGIC; 
  signal blk00000001_sig00000082 : STD_LOGIC; 
  signal blk00000001_sig00000081 : STD_LOGIC; 
  signal blk00000001_sig00000080 : STD_LOGIC; 
  signal blk00000001_sig0000007f : STD_LOGIC; 
  signal blk00000001_sig0000007e : STD_LOGIC; 
  signal blk00000001_sig0000007d : STD_LOGIC; 
  signal blk00000001_sig0000007c : STD_LOGIC; 
  signal blk00000001_sig0000007b : STD_LOGIC; 
  signal blk00000001_sig0000007a : STD_LOGIC; 
  signal blk00000001_sig00000079 : STD_LOGIC; 
  signal blk00000001_sig00000078 : STD_LOGIC; 
  signal blk00000001_sig00000077 : STD_LOGIC; 
  signal blk00000001_sig00000076 : STD_LOGIC; 
  signal blk00000001_sig00000075 : STD_LOGIC; 
  signal blk00000001_sig00000074 : STD_LOGIC; 
  signal blk00000001_sig00000073 : STD_LOGIC; 
  signal blk00000001_sig00000072 : STD_LOGIC; 
  signal blk00000001_sig00000071 : STD_LOGIC; 
  signal blk00000001_sig00000070 : STD_LOGIC; 
  signal blk00000001_sig0000006f : STD_LOGIC; 
  signal blk00000001_sig0000006e : STD_LOGIC; 
  signal blk00000001_sig0000006d : STD_LOGIC; 
  signal blk00000001_sig0000006c : STD_LOGIC; 
  signal blk00000001_sig0000006b : STD_LOGIC; 
  signal blk00000001_sig0000006a : STD_LOGIC; 
  signal blk00000001_sig00000069 : STD_LOGIC; 
  signal blk00000001_sig00000068 : STD_LOGIC; 
  signal blk00000001_sig00000067 : STD_LOGIC; 
  signal blk00000001_sig00000066 : STD_LOGIC; 
  signal blk00000001_sig00000065 : STD_LOGIC; 
  signal blk00000001_sig00000064 : STD_LOGIC; 
  signal blk00000001_sig00000063 : STD_LOGIC; 
  signal blk00000001_sig00000062 : STD_LOGIC; 
  signal blk00000001_sig00000061 : STD_LOGIC; 
  signal blk00000001_sig00000060 : STD_LOGIC; 
  signal blk00000001_sig0000005f : STD_LOGIC; 
  signal blk00000001_sig0000005e : STD_LOGIC; 
  signal blk00000001_blk00000022_sig00000201 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig00000200 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ff : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001fe : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001fd : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001fc : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001fb : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001fa : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f9 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f8 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f7 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f6 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f5 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f4 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f3 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f2 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f1 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001f0 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ef : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ee : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ed : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ec : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001eb : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001ea : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e9 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e8 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e7 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e6 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e5 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e4 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e3 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e2 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e1 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001e0 : STD_LOGIC; 
  signal blk00000001_blk00000022_sig000001df : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000282 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000281 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000280 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027f : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027e : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027d : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027c : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027b : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000027a : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000279 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000278 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000277 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000276 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000275 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000274 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000273 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000272 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000271 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000270 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026f : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026e : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026d : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026c : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026b : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000026a : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000269 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000268 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000267 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000266 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000265 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000264 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000263 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000262 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000261 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000260 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025f : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025e : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025d : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025c : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025b : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000025a : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000259 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000258 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000257 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000256 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000255 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000254 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000253 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000252 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000251 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig00000250 : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000024e : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000024d : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000024c : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000024b : STD_LOGIC; 
  signal blk00000001_blk000000ba_sig0000024a : STD_LOGIC; 
  signal blk00000001_blk00000117_sig000002a4 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig000002a3 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig000002a2 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig000002a1 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig000002a0 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029f : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029e : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029d : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029c : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029b : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000029a : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000299 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000298 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000297 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000296 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000295 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000294 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000293 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000292 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig00000291 : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000028e : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000028d : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000028c : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000028b : STD_LOGIC; 
  signal blk00000001_blk00000117_sig0000028a : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000033e : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000033d : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000033c : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000033b : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000033a : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000339 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000338 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000337 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000336 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000335 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000334 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000333 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000332 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000331 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000330 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032f : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032e : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032d : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032c : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032b : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000032a : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000329 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000328 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000327 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000326 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000325 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000324 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000323 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000322 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000321 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000320 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031f : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031e : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031d : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031c : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031b : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000031a : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000319 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000318 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000317 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000316 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000315 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000314 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000313 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000312 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000311 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000310 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030f : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030e : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030d : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030c : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030b : STD_LOGIC; 
  signal blk00000001_blk00000134_sig0000030a : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000309 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000308 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000307 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000306 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000305 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000304 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000303 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig00000302 : STD_LOGIC; 
  signal blk00000001_blk00000134_sig000002fe : STD_LOGIC; 
  signal blk00000001_blk00000134_sig000002fd : STD_LOGIC; 
  signal blk00000001_blk00000134_sig000002fc : STD_LOGIC; 
  signal blk00000001_blk00000134_sig000002fb : STD_LOGIC; 
  signal blk00000001_blk00000134_sig000002fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_sig00000754 : STD_LOGIC; 
  signal blk00000001_blk000001a2_sig00000753 : STD_LOGIC; 
  signal blk00000001_blk000001a2_sig00000592 : STD_LOGIC; 
  signal blk00000001_blk000001a2_sig0000053d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001402 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001401 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001400 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000013a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000139a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001399 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001398 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001397 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001396 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001395 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001394 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001393 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001392 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001391 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001390 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000138a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001389 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001388 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001387 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001386 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001385 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001384 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001383 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001382 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001381 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001380 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000137a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001379 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001378 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001377 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001376 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001375 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001374 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001373 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001372 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001371 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001370 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000136a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001369 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001368 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001367 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001366 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001365 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001364 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001363 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001362 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001361 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001360 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000135a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001359 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001358 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001357 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001356 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001355 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001354 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001353 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001352 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001351 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001350 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000134a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001349 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001348 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001347 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001346 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001345 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001344 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001343 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001342 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001341 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001340 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000133a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001339 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001338 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001337 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001336 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001335 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001334 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001333 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001332 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001331 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001330 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000132a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001329 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001328 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001327 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001326 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001325 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001324 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001323 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001322 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001321 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001320 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000131a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001319 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001318 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001317 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001316 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001315 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001314 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001313 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001312 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001311 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001310 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000130a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001309 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001308 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001307 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001306 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001305 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001304 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001303 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001302 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001301 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001300 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000012a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000129a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001299 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001298 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001297 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001296 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001295 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001294 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001293 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001292 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001291 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001290 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000128a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001289 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001288 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001287 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001286 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001285 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001284 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001283 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001282 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001281 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001280 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000127a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001279 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001278 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001277 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001276 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001275 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001274 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001273 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001272 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001271 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001270 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000126a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001269 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001268 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001267 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001266 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001265 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001264 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001263 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001262 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001261 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001260 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000125a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001259 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001258 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001257 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001256 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001255 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001254 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001253 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001252 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001251 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001250 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000124a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001249 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001248 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001247 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001246 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001245 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001244 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001243 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001242 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001241 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001240 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000123a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001239 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001238 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001237 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001236 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001235 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001234 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001233 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001232 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001231 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001230 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000122a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001229 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001228 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001227 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001226 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001225 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001224 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001223 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001222 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001221 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001220 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000121a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001219 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001218 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001217 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001216 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001215 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001214 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001213 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001212 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001211 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001210 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000120a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001209 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001208 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001207 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001206 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001205 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001204 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001203 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001202 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001201 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001200 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000011a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000119a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001199 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001198 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001197 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001196 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001195 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001194 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001193 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001192 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001191 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001190 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000118a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001189 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001188 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001187 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001186 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001185 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001184 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001183 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001182 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001181 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001180 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000117a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001179 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001178 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001177 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001176 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001175 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001174 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001173 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001172 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001171 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001170 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000116a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001169 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001168 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001167 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001166 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001165 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001164 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001163 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001162 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001161 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001160 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000115a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001159 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001158 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001157 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001156 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001155 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001154 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001153 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001152 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001151 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001150 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000114a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001149 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001148 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001147 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001146 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001145 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001144 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001143 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001142 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001141 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001140 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000113a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001139 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001138 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001137 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001136 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001135 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001134 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001133 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001132 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001131 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001130 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000112a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001129 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001128 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001127 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001126 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001125 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001124 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001123 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001122 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001121 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001120 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000111a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001119 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001118 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001117 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001116 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001115 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001114 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001113 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001112 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001111 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001110 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000110a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001109 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001108 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001107 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001106 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001105 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001104 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001103 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001102 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001101 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001100 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000010a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000109a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001099 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001098 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001097 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001096 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001095 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001094 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001093 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001092 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001091 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001090 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000108a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001089 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001088 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001087 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001086 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001085 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001084 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001083 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001082 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001081 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001080 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000107a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001079 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001078 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001077 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001076 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001075 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001074 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001073 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001072 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001071 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001070 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000106a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001069 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001068 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001067 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001066 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001065 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001064 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001063 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001062 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001061 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001060 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000105a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001059 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001058 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001057 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001056 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001055 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001054 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001053 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001052 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001051 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001050 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000104a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001049 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001048 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001047 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001046 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001045 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001044 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001043 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001042 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001041 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001040 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000103a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001039 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001038 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001037 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001036 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001035 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001034 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001033 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001032 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001031 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001030 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000102a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001029 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001028 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001027 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001026 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001025 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001024 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001023 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001022 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001021 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001020 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000101a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001019 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001018 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001017 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001016 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001015 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001014 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001013 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001012 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001011 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001010 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000100a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001009 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001008 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001007 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001006 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001005 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001004 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001003 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001002 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001001 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00001000 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ffe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ffd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ffc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ffb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ffa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ff0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000feb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fe0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fdf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fde : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fdd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fdc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fdb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fd0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fcf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fcd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fcc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fcb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fc0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fbf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fbe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fbd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fbc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fbb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000faf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000faa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000fa0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000f00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000efe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000efd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000efc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000efb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000efa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ef0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eeb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ee0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000edf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ede : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000edd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000edc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000edb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ed0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ecf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ece : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ecd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ecc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ecb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ec0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ebf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ebe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ebd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ebc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ebb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eaf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ead : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000eaa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ea0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000e00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dfe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dfd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dfc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dfb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dfa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000df0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000def : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ded : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000deb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000de0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ddf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dde : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ddd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ddc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ddb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dd0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dcf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dcd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dcc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dcb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dc0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dbf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dbe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dbd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dbc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dbb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000db0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000daf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000dab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000daa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000da0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000d00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cfe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cfd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cfc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cfb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cfa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cf0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ced : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ceb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ce0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cdf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cde : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cdd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cdc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cdb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cd0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ccf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ccd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ccc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ccb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cc0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cbf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cbe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cbd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cbc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cbb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000caf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000cab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000caa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ca0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000c00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bfe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bfd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bfc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bfb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bfa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bf0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000beb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000be0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bdf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bde : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bdd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bdc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bdb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bd0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bcf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bcd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bcc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bcb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bc0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bbf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bbe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bbd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bbc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bbb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000baf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000bab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000baa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ba0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000b00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000afe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000afd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000afc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000afb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000afa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000af0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aeb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ae0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000adf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ade : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000add : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000adc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000adb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ada : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ad0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000acf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ace : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000acd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000acc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000acb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ac0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000abf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000abe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000abd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000abc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000abb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000ab0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aaf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aaa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000aa0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a01 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000a00 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000009a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000099a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000999 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000998 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000997 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000996 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000995 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000994 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000993 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000992 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000991 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000990 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000098a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000989 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000988 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000987 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000986 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000985 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000984 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000983 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000982 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000981 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000980 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000097a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000979 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000978 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000977 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000976 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000975 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000974 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000973 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000972 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000971 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000970 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000096a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000969 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000968 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000967 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000966 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000965 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000964 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000963 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000962 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000961 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000960 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000095a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000959 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000958 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000957 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000956 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000955 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000954 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000953 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000952 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000951 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000950 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000094a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000949 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000948 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000947 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000946 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000945 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000944 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000943 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000942 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000941 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000940 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000093a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000939 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000938 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000937 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000936 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000935 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000934 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000933 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000932 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000931 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000930 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000092a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000929 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000928 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000927 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000926 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000925 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000924 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000923 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000922 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000921 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000920 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000091a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000919 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000918 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000917 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000916 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000915 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000914 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000913 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000912 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000911 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000910 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000090a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000909 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000908 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000907 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000906 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000905 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000904 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000903 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000902 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000901 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000900 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000008a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000089a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000899 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000898 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000897 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000896 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000895 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000894 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000893 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000892 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000891 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000890 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000088a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000889 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000888 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000887 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000886 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000885 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000884 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000883 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000882 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000881 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000880 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000087a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000879 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000878 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000877 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000876 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000875 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000874 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000873 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000872 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000871 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000870 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000086a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000869 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000868 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000867 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000866 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000865 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000864 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000863 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000862 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000861 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000860 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000085a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000859 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000858 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000857 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000856 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000855 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000854 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000853 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000852 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000851 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000850 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000084a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000849 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000848 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000847 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000846 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000845 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000844 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000843 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000842 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000841 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000840 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000083a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000839 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000838 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000837 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000836 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000835 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000834 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000833 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000832 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000831 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000830 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000082a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000829 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000828 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000827 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000826 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000825 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000824 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000823 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000822 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000821 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000820 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000081a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000819 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000818 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000817 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000816 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000815 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000814 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000813 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000812 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000811 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000810 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig0000080a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000809 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000808 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000807 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000806 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000805 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000804 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000803 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000802 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000801 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig00000800 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_sig000007c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001481 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001480 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001479 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001478 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001477 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001476 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001475 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001474 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001473 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001472 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001471 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001470 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001469 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001468 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001467 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001466 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001465 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001464 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001463 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001462 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001461 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001460 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001459 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001458 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001457 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001456 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001455 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001454 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001453 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001452 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001451 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001450 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001449 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001448 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001447 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001446 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001445 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001444 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001443 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig00001500 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001589 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001588 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001587 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001586 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001585 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001584 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001583 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001582 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001581 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001580 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001579 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001578 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001577 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001576 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001575 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001574 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001573 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001572 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001571 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001570 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001569 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001568 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001567 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001566 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001565 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001564 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001563 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001562 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001561 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001560 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001559 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001558 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001557 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001556 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001555 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001554 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001553 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001552 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001551 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001550 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001549 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001548 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001547 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001546 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001545 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001544 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001543 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001542 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001541 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001540 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000161a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001619 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001618 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001617 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001616 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001615 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001614 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001613 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001612 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001611 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001610 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001609 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001608 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001607 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001606 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001605 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001604 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001603 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001602 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001601 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001600 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001699 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001698 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001697 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001696 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001695 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001694 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001693 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001692 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001691 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001690 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001689 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001688 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001687 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001686 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001685 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001684 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001683 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001682 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001681 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001680 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001679 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001678 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001677 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001676 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001675 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001674 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001673 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001672 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001671 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001670 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001669 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001668 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001667 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001666 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001665 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001664 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001663 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001662 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001661 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001660 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001718 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001717 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001716 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001715 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001714 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001713 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001712 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001711 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001710 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001709 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001708 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001707 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001706 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001705 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001704 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001703 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001702 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001701 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001700 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016df : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016de : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016db : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016da : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001799 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001798 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001797 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001796 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001795 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001794 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001793 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001792 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001791 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001790 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001789 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001788 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001787 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001786 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001785 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001784 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001783 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001782 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001781 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001780 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001779 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001778 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001777 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001776 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001775 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001774 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001773 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001772 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001771 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001770 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001769 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001768 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001767 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001766 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001765 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001764 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001763 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001762 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001761 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001760 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001759 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001839 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001838 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001837 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001836 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001835 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001834 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001833 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001832 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001831 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001830 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001829 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001828 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001827 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001826 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001825 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001824 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001823 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001822 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001821 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001820 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001819 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001818 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001817 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001816 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001815 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001814 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001813 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001812 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001811 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001810 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001809 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001808 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001807 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001806 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001805 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001804 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001803 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001802 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001801 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001800 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ff : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ed : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017eb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001899 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001898 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001897 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001896 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001895 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001894 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001893 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001892 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001891 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001890 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001889 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001888 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001887 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001886 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001885 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001884 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001883 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001882 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001881 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001880 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000187f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001944 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001943 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001942 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001941 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001940 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001939 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001938 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001937 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001936 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001935 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001934 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001933 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001932 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001931 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001930 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001929 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001928 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001927 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001926 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001925 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001924 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001923 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001922 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001921 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001920 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001919 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001918 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001917 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001916 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001915 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001914 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001913 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001912 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001911 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001910 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001909 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001908 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001907 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001906 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001905 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001904 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001903 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019be : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019af : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019aa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001999 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001998 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001997 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001996 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001995 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001994 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001993 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001992 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001991 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001990 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001989 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001988 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001987 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ad0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ace : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a94 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a93 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a92 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a91 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a90 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a8f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bce : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bca : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbe : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c55 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c54 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c53 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c52 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c51 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c50 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c47 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c46 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c45 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c44 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c43 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c41 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c39 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c38 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c37 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c36 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c35 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c29 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c25 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cad : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d21 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d20 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d19 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d18 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d17 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d16 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d15 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d14 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d13 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d12 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d11 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d09 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d08 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d07 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d06 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d05 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d04 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d03 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d02 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d74 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d73 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d72 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d71 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001def : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dee : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ded : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dec : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001deb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dea : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dde : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddd : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e28 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e27 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e26 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e34 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e33 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e40 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e56 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e70 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e69 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e68 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e67 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e65 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e89 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e88 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e87 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e86 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e85 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e84 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e83 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e82 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e81 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e7f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e99 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e98 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e97 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e95 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eb0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaf : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eae : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ead : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eac : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eab : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001ebb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eba : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eb9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec7 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec3 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec2 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001edb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001eda : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee6 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee5 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee4 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef1 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef0 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001eef : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efc : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efb : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efa : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f10 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f24 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f23 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f32 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f2f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f4a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f49 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f48 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f64 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f63 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f62 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f61 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f60 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5f : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f59 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f58 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f57 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7e : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7d : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7c : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7b : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7a : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f79 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f78 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f77 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f76 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f75 : STD_LOGIC; 
  signal blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f74 : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000043_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000042_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000041_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000040_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk0000003a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000039_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000038_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000022_blk00000037_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk0000010c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk0000010b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk00000101_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk00000100_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ff_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000fe_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000fd_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000fc_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000fb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000fa_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f2_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000f0_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ef_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ee_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ed_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ec_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000eb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000ea_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e8_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e6_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e4_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000000ba_blk000000e3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000117_blk00000122_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000166_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000165_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000164_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000163_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000162_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000161_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000160_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000015a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000159_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000158_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000157_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000156_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000155_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000154_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000153_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000152_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000151_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000150_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014d_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014c_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk0000014a_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000149_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000148_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000147_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000146_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000145_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000144_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000143_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000142_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000141_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000137_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk00000134_blk00000136_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_43_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_42_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_41_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_40_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_39_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_38_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_37_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_36_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_35_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_34_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_33_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_32_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PATTERNBDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_MULTSIGNOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYCASCOUT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_UNDERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PATTERNDETECT_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_OVERFLOW_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_28_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_27_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_26_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_25_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_24_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_23_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_22_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_21_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_20_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_19_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_18_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_17_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_16_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_47_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_46_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_45_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_44_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000115b_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001159_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001157_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001155_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001153_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_14_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_13_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_12_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_11_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_10_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_9_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_8_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_7_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_6_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_5_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_4_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_2_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIPBDIP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIPBDIP_0_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DOPADOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DOPBDOP_1_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fce_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fcd_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fc2_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fc0_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fb4_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000fb2_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f86_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f84_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f80_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f7e_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f10_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000056d_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000056c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000056b_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000056a_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000569_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000568_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000053b_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000053a_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000539_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000538_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000537_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000536_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000509_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000508_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000507_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000506_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000505_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000504_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d7_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d6_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d5_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d4_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004d2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a5_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a4_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a3_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a2_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a1_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk000004a0_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000473_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000472_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000471_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000470_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000046f_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000046e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000441_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000440_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000043f_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000043e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000043d_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000043c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040f_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040e_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040d_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040c_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040b_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk0000040a_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c4f_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DOP_3_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_30_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_29_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000de1_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de7_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000ded_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df3_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000df9_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000ed9_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000edf_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee5_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000eeb_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000ef1_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef7_Q31_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f19_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f18_Q_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1e_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f25_Q15_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f54_O_UNCONNECTED : STD_LOGIC; 
begin
  m_axis_data_tuser(15) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(14) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(13) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(12) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(11) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(10) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(9) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(8) <= NlwRenamedSig_OI_m_axis_data_tuser_8_Q;
  m_axis_data_tuser(7) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_data_tuser(6) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(7) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(6) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(5) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(4) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(3) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(2) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  m_axis_status_tdata(1) <= NlwRenamedSig_OI_m_axis_data_tuser_10_Q;
  s_axis_config_tready <= NlwRenamedSig_OI_s_axis_config_tready;
  s_axis_data_tready <= NlwRenamedSig_OI_s_axis_data_tready;
  m_axis_data_tvalid <= NlwRenamedSig_OI_m_axis_data_tvalid;
  m_axis_status_tvalid <= NlwRenamedSig_OI_m_axis_status_tvalid;
  event_frame_started <= NlwRenamedSig_OI_event_frame_started;
  event_tlast_missing <= NlwRenamedSig_OI_event_tlast_missing;
  event_fft_overflow <= NlwRenamedSig_OI_event_fft_overflow;
  event_status_channel_halt <= NlwRenamedSig_OI_event_status_channel_halt;
  event_data_in_channel_halt <= NlwRenamedSig_OI_event_data_in_channel_halt;
  event_data_out_channel_halt <= NlwRenamedSig_OI_event_data_out_channel_halt;
  blk00000001_blk000011da : LUT6
    generic map(
      INIT => X"FFFFFFFF44404040"
    )
    port map (
      I0 => blk00000001_sig000000ce,
      I1 => blk00000001_sig000000e8,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig000000d0,
      I4 => blk00000001_sig000000e7,
      I5 => blk00000001_sig000001ba,
      O => blk00000001_sig000001be
    );
  blk00000001_blk000011d9 : LUT5
    generic map(
      INIT => X"88888000"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig000001bb,
      I2 => blk00000001_sig000000e7,
      I3 => blk00000001_sig000000d0,
      I4 => blk00000001_sig000000c7,
      O => blk00000001_sig000001bd
    );
  blk00000001_blk000011d8 : MUXF7
    port map (
      I0 => blk00000001_sig000001bd,
      I1 => blk00000001_sig000001be,
      S => NlwRenamedSig_OI_event_frame_started,
      O => blk00000001_sig000001ae
    );
  blk00000001_blk000011d7 : INV
    port map (
      I => aresetn,
      O => blk00000001_sig000000d7
    );
  blk00000001_blk000011d6 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig000000cf,
      I1 => blk00000001_sig000001bc,
      I2 => blk00000001_sig000000f4,
      O => blk00000001_sig000001b4
    );
  blk00000001_blk000011d5 : LUT6
    generic map(
      INIT => X"DF8A8A8A8A8A8A8A"
    )
    port map (
      I0 => blk00000001_sig000000eb,
      I1 => blk00000001_sig000000fd,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_sig000000cf,
      I4 => blk00000001_sig000000c9,
      I5 => blk00000001_sig000000d1,
      O => blk00000001_sig000001ac
    );
  blk00000001_blk000011d4 : LUT6
    generic map(
      INIT => X"00020002FFFF0002"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig000000ff,
      I2 => blk00000001_sig000000f1,
      I3 => blk00000001_sig000000d0,
      I4 => NlwRenamedSig_OI_event_tlast_missing,
      I5 => aclken,
      O => blk00000001_sig000001ad
    );
  blk00000001_blk000011d3 : LUT5
    generic map(
      INIT => X"444444E4"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_event_data_in_channel_halt,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig000000f1,
      I4 => blk00000001_sig000000fe,
      O => blk00000001_sig000001b2
    );
  blk00000001_blk000011d2 : LUT6
    generic map(
      INIT => X"FFFFFFFF02000000"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig000000fe,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig000000e8,
      I4 => blk00000001_sig000000e6,
      I5 => blk00000001_sig000000f1,
      O => blk00000001_sig000001af
    );
  blk00000001_blk000011d1 : LUT4
    generic map(
      INIT => X"BA10"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => blk00000001_sig00000097,
      I2 => blk00000001_sig000000fa,
      I3 => blk00000001_sig000000f5,
      O => blk00000001_sig000001b3
    );
  blk00000001_blk000011d0 : LUT5
    generic map(
      INIT => X"04550400"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => blk00000001_sig000000c9,
      I2 => blk00000001_sig000000ca,
      I3 => blk00000001_sig0000009a,
      I4 => blk00000001_sig000000f2,
      O => blk00000001_sig000001b8
    );
  blk00000001_blk000011cf : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => aclken,
      I2 => blk00000001_sig000000fc,
      I3 => blk00000001_sig000000c9,
      I4 => NlwRenamedSig_OI_event_data_out_channel_halt,
      O => blk00000001_sig000001b7
    );
  blk00000001_blk000011ce : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => aclken,
      I2 => blk00000001_sig000000eb,
      I3 => blk00000001_sig000000fd,
      I4 => NlwRenamedSig_OI_event_status_channel_halt,
      O => blk00000001_sig000001b6
    );
  blk00000001_blk000011cd : LUT6
    generic map(
      INIT => X"5410101010101010"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_event_fft_overflow,
      I3 => m_axis_data_tready,
      I4 => NlwRenamedSig_OI_m_axis_data_tuser_8_Q,
      I5 => NlwRenamedSig_OI_m_axis_data_tvalid,
      O => blk00000001_sig000001b5
    );
  blk00000001_blk000011cc : LUT6
    generic map(
      INIT => X"AAAAAAEAAAAAAA2A"
    )
    port map (
      I0 => blk00000001_sig000000f4,
      I1 => blk00000001_sig000000d1,
      I2 => blk00000001_sig000000c9,
      I3 => blk00000001_sig000000f6,
      I4 => blk00000001_sig000000eb,
      I5 => blk00000001_sig000000cb,
      O => blk00000001_sig000001bc
    );
  blk00000001_blk000011cb : LUT6
    generic map(
      INIT => X"FFFFFFFFAAAAAA6A"
    )
    port map (
      I0 => blk00000001_sig000000d1,
      I1 => blk00000001_sig000000c9,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_sig000000ca,
      I4 => blk00000001_sig000000f6,
      I5 => blk00000001_sig000000e0,
      O => blk00000001_sig000001ab
    );
  blk00000001_blk000011ca : LUT4
    generic map(
      INIT => X"F888"
    )
    port map (
      I0 => blk00000001_sig000000e7,
      I1 => blk00000001_sig000000d0,
      I2 => blk00000001_sig000000e8,
      I3 => blk00000001_sig000000c7,
      O => blk00000001_sig000000de
    );
  blk00000001_blk000011c9 : LUT6
    generic map(
      INIT => X"2020200020002000"
    )
    port map (
      I0 => blk00000001_sig000000e8,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000f3,
      I3 => blk00000001_sig000000c7,
      I4 => blk00000001_sig000000e7,
      I5 => blk00000001_sig000000d0,
      O => blk00000001_sig000000df
    );
  blk00000001_blk000011c8 : LUT5
    generic map(
      INIT => X"0040AAEA"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig000000fe,
      I2 => blk00000001_sig00000159,
      I3 => blk00000001_sig000000e4,
      I4 => blk00000001_sig00000113,
      O => blk00000001_sig000001b1
    );
  blk00000001_blk000011c7 : LUT4
    generic map(
      INIT => X"FFA6"
    )
    port map (
      I0 => blk00000001_sig000000ec,
      I1 => blk00000001_sig000000d6,
      I2 => blk00000001_sig000000d1,
      I3 => blk00000001_sig000000e0,
      O => blk00000001_sig000001aa
    );
  blk00000001_blk000011c6 : LUT5
    generic map(
      INIT => X"FFFFAA9A"
    )
    port map (
      I0 => blk00000001_sig000000ed,
      I1 => blk00000001_sig000000d1,
      I2 => blk00000001_sig000000d6,
      I3 => blk00000001_sig000000ec,
      I4 => blk00000001_sig000000e0,
      O => blk00000001_sig000001a9
    );
  blk00000001_blk000011c5 : LUT6
    generic map(
      INIT => X"FFFFFFFFAAAAA9AA"
    )
    port map (
      I0 => blk00000001_sig000000ee,
      I1 => blk00000001_sig000000d1,
      I2 => blk00000001_sig000000ec,
      I3 => blk00000001_sig000000d6,
      I4 => blk00000001_sig000000ed,
      I5 => blk00000001_sig000000e0,
      O => blk00000001_sig000001a8
    );
  blk00000001_blk000011c4 : LUT6
    generic map(
      INIT => X"FFFFFFFFAA8AAAAA"
    )
    port map (
      I0 => blk00000001_sig000000fe,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig000000f6,
      I4 => blk00000001_sig0000009a,
      I5 => blk00000001_sig00000112,
      O => blk00000001_sig000001b0
    );
  blk00000001_blk000011c3 : LUT4
    generic map(
      INIT => X"DFFF"
    )
    port map (
      I0 => blk00000001_sig000000c7,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000ff,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_sig000001b9
    );
  blk00000001_blk000011c2 : LUT6
    generic map(
      INIT => X"00002000AAAAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      I4 => blk00000001_sig000000f6,
      I5 => blk00000001_sig000000fe,
      O => blk00000001_sig00000113
    );
  blk00000001_blk000011c1 : LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      I0 => blk00000001_sig000000ca,
      I1 => blk00000001_sig000000c9,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_sig000000f6,
      O => blk00000001_sig000000d6
    );
  blk00000001_blk000011c0 : LUT2
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_sig000000e8,
      I1 => blk00000001_sig000000f1,
      O => blk00000001_sig000001bb
    );
  blk00000001_blk000011bf : LUT6
    generic map(
      INIT => X"555555554A4AAA4A"
    )
    port map (
      I0 => blk00000001_sig000000f8,
      I1 => blk00000001_sig000000f9,
      I2 => aclken,
      I3 => blk00000001_sig000000d0,
      I4 => blk00000001_sig000001b9,
      I5 => blk00000001_sig000000cd,
      O => blk00000001_sig000000d3
    );
  blk00000001_blk000011be : LUT6
    generic map(
      INIT => X"77777777AEAEEEAE"
    )
    port map (
      I0 => blk00000001_sig000000f9,
      I1 => blk00000001_sig000000f8,
      I2 => aclken,
      I3 => blk00000001_sig000000d0,
      I4 => blk00000001_sig000001b9,
      I5 => blk00000001_sig000000cd,
      O => blk00000001_sig000000d8
    );
  blk00000001_blk000011bd : LUT6
    generic map(
      INIT => X"3C3C3C3CD0F0D0D0"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000f8,
      I2 => blk00000001_sig000000f9,
      I3 => blk00000001_sig000001b9,
      I4 => blk00000001_sig000000d0,
      I5 => blk00000001_sig000000cd,
      O => blk00000001_sig000000d2
    );
  blk00000001_blk000011bc : LUT6
    generic map(
      INIT => X"AAAAAAAAAAAAAAA9"
    )
    port map (
      I0 => blk00000001_sig000000f0,
      I1 => blk00000001_sig000000ef,
      I2 => blk00000001_sig000000ee,
      I3 => blk00000001_sig000000ed,
      I4 => blk00000001_sig000000ec,
      I5 => blk00000001_sig000000d1,
      O => blk00000001_sig000000d4
    );
  blk00000001_blk000011bb : LUT4
    generic map(
      INIT => X"FFD8"
    )
    port map (
      I0 => blk00000001_sig000000d6,
      I1 => blk00000001_sig000000d5,
      I2 => blk00000001_sig000000ef,
      I3 => blk00000001_sig000000e0,
      O => blk00000001_sig000001a7
    );
  blk00000001_blk000011ba : LUT4
    generic map(
      INIT => X"FFD8"
    )
    port map (
      I0 => blk00000001_sig000000d6,
      I1 => blk00000001_sig000000d4,
      I2 => blk00000001_sig000000f0,
      I3 => blk00000001_sig000000e0,
      O => blk00000001_sig000001a6
    );
  blk00000001_blk000011b9 : LUT2
    generic map(
      INIT => X"7"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_event_frame_started,
      O => blk00000001_sig000001ba
    );
  blk00000001_blk000011b8 : LUT5
    generic map(
      INIT => X"55557555"
    )
    port map (
      I0 => blk00000001_sig000000fe,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      I4 => blk00000001_sig000000f6,
      O => blk00000001_sig00000136
    );
  blk00000001_blk000011b7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b8,
      Q => blk00000001_sig000000f2
    );
  blk00000001_blk000011b6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b7,
      Q => NlwRenamedSig_OI_event_data_out_channel_halt
    );
  blk00000001_blk000011b5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b6,
      Q => NlwRenamedSig_OI_event_status_channel_halt
    );
  blk00000001_blk000011b4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b5,
      Q => NlwRenamedSig_OI_event_fft_overflow
    );
  blk00000001_blk000011b3 : FD
    port map (
      C => aclk,
      D => blk00000001_sig000001b4,
      Q => blk00000001_sig000000f4
    );
  blk00000001_blk000011b2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b3,
      Q => blk00000001_sig000000f5
    );
  blk00000001_blk000011b1 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b2,
      R => blk00000001_sig000000f6,
      Q => NlwRenamedSig_OI_event_data_in_channel_halt
    );
  blk00000001_blk000011b0 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b1,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000137
    );
  blk00000001_blk000011af : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001b0,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000fe
    );
  blk00000001_blk000011ae : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001af,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000f1
    );
  blk00000001_blk000011ad : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001ae,
      R => blk00000001_sig000000f6,
      Q => NlwRenamedSig_OI_event_frame_started
    );
  blk00000001_blk000011ac : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001ad,
      R => blk00000001_sig000000f6,
      Q => NlwRenamedSig_OI_event_tlast_missing
    );
  blk00000001_blk000011ab : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001ac,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000eb
    );
  blk00000001_blk000011aa : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001ab,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000d1
    );
  blk00000001_blk000011a9 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001aa,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ec
    );
  blk00000001_blk000011a8 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001a9,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ed
    );
  blk00000001_blk000011a7 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001a8,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ee
    );
  blk00000001_blk000011a6 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001a7,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ef
    );
  blk00000001_blk000011a5 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000001a6,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000f0
    );
  blk00000001_blk000011a4 : LUT6
    generic map(
      INIT => X"C8C8C0C800000000"
    )
    port map (
      I0 => blk00000001_sig000000fe,
      I1 => blk00000001_sig000001a4,
      I2 => blk00000001_sig000001a2,
      I3 => blk00000001_sig000000d0,
      I4 => blk00000001_sig000001a5,
      I5 => blk00000001_sig000001a3,
      O => blk00000001_sig000000da
    );
  blk00000001_blk000011a3 : LUT5
    generic map(
      INIT => X"FF8FFFAF"
    )
    port map (
      I0 => blk00000001_sig0000015a,
      I1 => blk00000001_sig00000159,
      I2 => blk00000001_sig000000fe,
      I3 => blk00000001_sig00000137,
      I4 => blk00000001_sig000000e4,
      O => blk00000001_sig000001a5
    );
  blk00000001_blk000011a2 : LUT3
    generic map(
      INIT => X"2A"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000fd,
      I2 => blk00000001_sig000000eb,
      O => blk00000001_sig000001a4
    );
  blk00000001_blk000011a1 : LUT6
    generic map(
      INIT => X"13111F1F11111F1F"
    )
    port map (
      I0 => blk00000001_sig000000fb,
      I1 => blk00000001_sig000000fc,
      I2 => blk00000001_sig000000c8,
      I3 => blk00000001_sig000000d1,
      I4 => blk00000001_sig000000c9,
      I5 => blk00000001_sig000000cf,
      O => blk00000001_sig000001a3
    );
  blk00000001_blk000011a0 : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => blk00000001_sig000000f1,
      I1 => blk00000001_sig000000c7,
      O => blk00000001_sig000001a2
    );
  blk00000001_blk0000119f : LUT6
    generic map(
      INIT => X"0000200000000000"
    )
    port map (
      I0 => blk00000001_sig000000ff,
      I1 => blk00000001_sig000000f1,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      I4 => blk00000001_sig000001a1,
      I5 => blk00000001_sig000000d0,
      O => blk00000001_sig000000cd
    );
  blk00000001_blk0000119e : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig000000f9,
      I2 => blk00000001_sig000000f8,
      O => blk00000001_sig000001a1
    );
  blk00000001_blk0000119d : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => NlwRenamedSig_OI_s_axis_data_tready,
      I1 => aclken,
      I2 => blk00000001_sig000000f6,
      I3 => s_axis_data_tvalid,
      O => blk00000001_sig0000017d
    );
  blk00000001_blk0000119c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig0000017f,
      I2 => NlwRenamedSig_OI_s_axis_data_tready,
      O => blk00000001_sig0000017c
    );
  blk00000001_blk0000119b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000141,
      I2 => blk00000001_sig00000164,
      O => blk00000001_sig0000011e
    );
  blk00000001_blk0000119a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000140,
      I2 => blk00000001_sig00000163,
      O => blk00000001_sig0000011d
    );
  blk00000001_blk00001199 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013f,
      I2 => blk00000001_sig00000162,
      O => blk00000001_sig0000011c
    );
  blk00000001_blk00001198 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013e,
      I2 => blk00000001_sig00000161,
      O => blk00000001_sig0000011b
    );
  blk00000001_blk00001197 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013d,
      I2 => blk00000001_sig00000160,
      O => blk00000001_sig0000011a
    );
  blk00000001_blk00001196 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013c,
      I2 => blk00000001_sig0000015f,
      O => blk00000001_sig00000119
    );
  blk00000001_blk00001195 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000158,
      I2 => blk00000001_sig0000017b,
      O => blk00000001_sig00000135
    );
  blk00000001_blk00001194 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000157,
      I2 => blk00000001_sig0000017a,
      O => blk00000001_sig00000134
    );
  blk00000001_blk00001193 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000156,
      I2 => blk00000001_sig00000179,
      O => blk00000001_sig00000133
    );
  blk00000001_blk00001192 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013b,
      I2 => blk00000001_sig0000015e,
      O => blk00000001_sig00000118
    );
  blk00000001_blk00001191 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000155,
      I2 => blk00000001_sig00000178,
      O => blk00000001_sig00000132
    );
  blk00000001_blk00001190 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000154,
      I2 => blk00000001_sig00000177,
      O => blk00000001_sig00000131
    );
  blk00000001_blk0000118f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000153,
      I2 => blk00000001_sig00000176,
      O => blk00000001_sig00000130
    );
  blk00000001_blk0000118e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000152,
      I2 => blk00000001_sig00000175,
      O => blk00000001_sig0000012f
    );
  blk00000001_blk0000118d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000151,
      I2 => blk00000001_sig00000174,
      O => blk00000001_sig0000012e
    );
  blk00000001_blk0000118c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000150,
      I2 => blk00000001_sig00000173,
      O => blk00000001_sig0000012d
    );
  blk00000001_blk0000118b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014f,
      I2 => blk00000001_sig00000172,
      O => blk00000001_sig0000012c
    );
  blk00000001_blk0000118a : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014e,
      I2 => blk00000001_sig00000171,
      O => blk00000001_sig0000012b
    );
  blk00000001_blk00001189 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014d,
      I2 => blk00000001_sig00000170,
      O => blk00000001_sig0000012a
    );
  blk00000001_blk00001188 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014c,
      I2 => blk00000001_sig0000016f,
      O => blk00000001_sig00000129
    );
  blk00000001_blk00001187 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000013a,
      I2 => blk00000001_sig0000015d,
      O => blk00000001_sig00000117
    );
  blk00000001_blk00001186 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014b,
      I2 => blk00000001_sig0000016e,
      O => blk00000001_sig00000128
    );
  blk00000001_blk00001185 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig0000014a,
      I2 => blk00000001_sig0000016d,
      O => blk00000001_sig00000127
    );
  blk00000001_blk00001184 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000149,
      I2 => blk00000001_sig0000016c,
      O => blk00000001_sig00000126
    );
  blk00000001_blk00001183 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000148,
      I2 => blk00000001_sig0000016b,
      O => blk00000001_sig00000125
    );
  blk00000001_blk00001182 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000147,
      I2 => blk00000001_sig0000016a,
      O => blk00000001_sig00000124
    );
  blk00000001_blk00001181 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000146,
      I2 => blk00000001_sig00000169,
      O => blk00000001_sig00000123
    );
  blk00000001_blk00001180 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000145,
      I2 => blk00000001_sig00000168,
      O => blk00000001_sig00000122
    );
  blk00000001_blk0000117f : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000144,
      I2 => blk00000001_sig00000167,
      O => blk00000001_sig00000121
    );
  blk00000001_blk0000117e : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000143,
      I2 => blk00000001_sig00000166,
      O => blk00000001_sig00000120
    );
  blk00000001_blk0000117d : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000142,
      I2 => blk00000001_sig00000165,
      O => blk00000001_sig0000011f
    );
  blk00000001_blk0000117c : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000139,
      I2 => blk00000001_sig0000015c,
      O => blk00000001_sig00000116
    );
  blk00000001_blk0000117b : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000138,
      I2 => blk00000001_sig0000015b,
      O => blk00000001_sig00000115
    );
  blk00000001_blk0000117a : LUT4
    generic map(
      INIT => X"0040"
    )
    port map (
      I0 => blk00000001_sig00000137,
      I1 => blk00000001_sig00000159,
      I2 => blk00000001_sig000000fe,
      I3 => blk00000001_sig000000e4,
      O => blk00000001_sig00000114
    );
  blk00000001_blk00001179 : LUT4
    generic map(
      INIT => X"FA32"
    )
    port map (
      I0 => blk00000001_sig00000159,
      I1 => blk00000001_sig000000fe,
      I2 => blk00000001_sig00000137,
      I3 => blk00000001_sig000000e4,
      O => blk00000001_sig00000112
    );
  blk00000001_blk00001178 : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => NlwRenamedSig_OI_s_axis_config_tready,
      I1 => aclken,
      I2 => blk00000001_sig000000f6,
      I3 => s_axis_config_tvalid,
      O => blk00000001_sig00000102
    );
  blk00000001_blk00001177 : LUT3
    generic map(
      INIT => X"D8"
    )
    port map (
      I0 => aclken,
      I1 => blk00000001_sig00000104,
      I2 => NlwRenamedSig_OI_s_axis_config_tready,
      O => blk00000001_sig00000101
    );
  blk00000001_blk00001176 : LUT4
    generic map(
      INIT => X"F222"
    )
    port map (
      I0 => blk00000001_sig000000e5,
      I1 => blk00000001_sig000000c9,
      I2 => blk00000001_sig000000e6,
      I3 => blk00000001_sig000000c8,
      O => blk00000001_sig000000dd
    );
  blk00000001_blk00001175 : LUT4
    generic map(
      INIT => X"A0EC"
    )
    port map (
      I0 => blk00000001_sig000000ea,
      I1 => blk00000001_sig000000e8,
      I2 => blk00000001_sig000000fe,
      I3 => blk00000001_sig000000c7,
      O => blk00000001_sig00000096
    );
  blk00000001_blk00001174 : LUT4
    generic map(
      INIT => X"22F2"
    )
    port map (
      I0 => blk00000001_sig000000ea,
      I1 => blk00000001_sig000000fe,
      I2 => blk00000001_sig000000e9,
      I3 => blk00000001_sig000000c9,
      O => blk00000001_sig000000db
    );
  blk00000001_blk00001173 : LUT6
    generic map(
      INIT => X"7FFFFFFFFFFFFFFF"
    )
    port map (
      I0 => blk00000001_sig0000009e,
      I1 => blk00000001_sig0000009d,
      I2 => blk00000001_sig0000009c,
      I3 => blk00000001_sig0000009b,
      I4 => blk00000001_sig000000a0,
      I5 => blk00000001_sig0000009f,
      O => blk00000001_sig000000d0
    );
  blk00000001_blk00001172 : LUT5
    generic map(
      INIT => X"0202FF02"
    )
    port map (
      I0 => blk00000001_sig000000e7,
      I1 => blk00000001_sig000000d0,
      I2 => blk00000001_sig000000f1,
      I3 => blk00000001_sig000000e6,
      I4 => blk00000001_sig000000c8,
      O => blk00000001_sig000000d9
    );
  blk00000001_blk00001171 : LUT5
    generic map(
      INIT => X"00000001"
    )
    port map (
      I0 => blk00000001_sig000000ec,
      I1 => blk00000001_sig000000ed,
      I2 => blk00000001_sig000000ee,
      I3 => blk00000001_sig000000ef,
      I4 => blk00000001_sig000000f0,
      O => blk00000001_sig000000cf
    );
  blk00000001_blk00001170 : LUT2
    generic map(
      INIT => X"B"
    )
    port map (
      I0 => blk00000001_sig000000f1,
      I1 => blk00000001_sig0000009a,
      O => blk00000001_sig000000ce
    );
  blk00000001_blk0000116f : LUT3
    generic map(
      INIT => X"20"
    )
    port map (
      I0 => blk00000001_sig000000c9,
      I1 => blk00000001_sig000000f6,
      I2 => blk00000001_sig0000009a,
      O => blk00000001_sig000000e2
    );
  blk00000001_blk0000116e : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig000000c9,
      I1 => blk00000001_sig000000d1,
      I2 => blk00000001_sig000000cf,
      O => blk00000001_sig000000e3
    );
  blk00000001_blk0000116d : LUT6
    generic map(
      INIT => X"0020AAAA00200020"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig000000f2,
      I2 => blk00000001_sig000000c9,
      I3 => blk00000001_sig000000ca,
      I4 => blk00000001_sig000000d1,
      I5 => blk00000001_sig000000cf,
      O => blk00000001_sig000000e0
    );
  blk00000001_blk0000116c : LUT3
    generic map(
      INIT => X"A8"
    )
    port map (
      I0 => blk00000001_sig000000c9,
      I1 => blk00000001_sig000000e5,
      I2 => blk00000001_sig000000e9,
      O => blk00000001_sig000000dc
    );
  blk00000001_blk0000116b : LUT4
    generic map(
      INIT => X"0400"
    )
    port map (
      I0 => blk00000001_sig000000f1,
      I1 => blk00000001_sig000000c7,
      I2 => blk00000001_sig000000f6,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_sig000000e4
    );
  blk00000001_blk0000116a : LUT3
    generic map(
      INIT => X"40"
    )
    port map (
      I0 => blk00000001_sig000000fd,
      I1 => blk00000001_sig000000eb,
      I2 => blk00000001_sig0000009a,
      O => blk00000001_sig000000e1
    );
  blk00000001_blk00001169 : LUT5
    generic map(
      INIT => X"AAAAAAA9"
    )
    port map (
      I0 => blk00000001_sig000000ef,
      I1 => blk00000001_sig000000d1,
      I2 => blk00000001_sig000000ec,
      I3 => blk00000001_sig000000ed,
      I4 => blk00000001_sig000000ee,
      O => blk00000001_sig000000d5
    );
  blk00000001_blk000000b9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tlast,
      Q => blk00000001_sig00000180
    );
  blk00000001_blk000000b8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(0),
      Q => blk00000001_sig00000181
    );
  blk00000001_blk000000b7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(1),
      Q => blk00000001_sig00000182
    );
  blk00000001_blk000000b6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(2),
      Q => blk00000001_sig00000183
    );
  blk00000001_blk000000b5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(3),
      Q => blk00000001_sig00000184
    );
  blk00000001_blk000000b4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(4),
      Q => blk00000001_sig00000185
    );
  blk00000001_blk000000b3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(5),
      Q => blk00000001_sig00000186
    );
  blk00000001_blk000000b2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(6),
      Q => blk00000001_sig00000187
    );
  blk00000001_blk000000b1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(7),
      Q => blk00000001_sig00000188
    );
  blk00000001_blk000000b0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(8),
      Q => blk00000001_sig00000189
    );
  blk00000001_blk000000af : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(9),
      Q => blk00000001_sig0000018a
    );
  blk00000001_blk000000ae : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(10),
      Q => blk00000001_sig0000018b
    );
  blk00000001_blk000000ad : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(11),
      Q => blk00000001_sig0000018c
    );
  blk00000001_blk000000ac : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(12),
      Q => blk00000001_sig0000018d
    );
  blk00000001_blk000000ab : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(13),
      Q => blk00000001_sig0000018e
    );
  blk00000001_blk000000aa : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(14),
      Q => blk00000001_sig0000018f
    );
  blk00000001_blk000000a9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(15),
      Q => blk00000001_sig00000190
    );
  blk00000001_blk000000a8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(16),
      Q => blk00000001_sig00000191
    );
  blk00000001_blk000000a7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(17),
      Q => blk00000001_sig00000192
    );
  blk00000001_blk000000a6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(18),
      Q => blk00000001_sig00000193
    );
  blk00000001_blk000000a5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(19),
      Q => blk00000001_sig00000194
    );
  blk00000001_blk000000a4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(20),
      Q => blk00000001_sig00000195
    );
  blk00000001_blk000000a3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(21),
      Q => blk00000001_sig00000196
    );
  blk00000001_blk000000a2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(22),
      Q => blk00000001_sig00000197
    );
  blk00000001_blk000000a1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(23),
      Q => blk00000001_sig00000198
    );
  blk00000001_blk000000a0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(24),
      Q => blk00000001_sig00000199
    );
  blk00000001_blk0000009f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(25),
      Q => blk00000001_sig0000019a
    );
  blk00000001_blk0000009e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(26),
      Q => blk00000001_sig0000019b
    );
  blk00000001_blk0000009d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(27),
      Q => blk00000001_sig0000019c
    );
  blk00000001_blk0000009c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(28),
      Q => blk00000001_sig0000019d
    );
  blk00000001_blk0000009b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(29),
      Q => blk00000001_sig0000019e
    );
  blk00000001_blk0000009a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(30),
      Q => blk00000001_sig0000019f
    );
  blk00000001_blk00000099 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_data_tdata(31),
      Q => blk00000001_sig000001a0
    );
  blk00000001_blk00000098 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig0000017c,
      Q => NlwRenamedSig_OI_s_axis_data_tready
    );
  blk00000001_blk00000097 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig0000017d,
      Q => blk00000001_sig0000017e
    );
  blk00000001_blk00000096 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000015b,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000138
    );
  blk00000001_blk00000095 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000015c,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000139
    );
  blk00000001_blk00000094 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000015d,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013a
    );
  blk00000001_blk00000093 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000015e,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013b
    );
  blk00000001_blk00000092 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000015f,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013c
    );
  blk00000001_blk00000091 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000160,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013d
    );
  blk00000001_blk00000090 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000161,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013e
    );
  blk00000001_blk0000008f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000162,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000013f
    );
  blk00000001_blk0000008e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000163,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000140
    );
  blk00000001_blk0000008d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000164,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000141
    );
  blk00000001_blk0000008c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000165,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000142
    );
  blk00000001_blk0000008b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000166,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000143
    );
  blk00000001_blk0000008a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000167,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000144
    );
  blk00000001_blk00000089 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000168,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000145
    );
  blk00000001_blk00000088 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000169,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000146
    );
  blk00000001_blk00000087 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016a,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000147
    );
  blk00000001_blk00000086 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016b,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000148
    );
  blk00000001_blk00000085 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016c,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000149
    );
  blk00000001_blk00000084 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016d,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014a
    );
  blk00000001_blk00000083 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016e,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014b
    );
  blk00000001_blk00000082 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000016f,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014c
    );
  blk00000001_blk00000081 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000170,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014d
    );
  blk00000001_blk00000080 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000171,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014e
    );
  blk00000001_blk0000007f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000172,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000014f
    );
  blk00000001_blk0000007e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000173,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000150
    );
  blk00000001_blk0000007d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000174,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000151
    );
  blk00000001_blk0000007c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000175,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000152
    );
  blk00000001_blk0000007b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000176,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000153
    );
  blk00000001_blk0000007a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000177,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000154
    );
  blk00000001_blk00000079 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000178,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000155
    );
  blk00000001_blk00000078 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig00000179,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000156
    );
  blk00000001_blk00000077 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000017a,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000157
    );
  blk00000001_blk00000076 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000114,
      D => blk00000001_sig0000017b,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000158
    );
  blk00000001_blk00000075 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000115,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ff
    );
  blk00000001_blk00000074 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000116,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000073
    );
  blk00000001_blk00000073 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000117,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000072
    );
  blk00000001_blk00000072 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000118,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000071
    );
  blk00000001_blk00000071 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000119,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000070
    );
  blk00000001_blk00000070 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011a,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006f
    );
  blk00000001_blk0000006f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011b,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006e
    );
  blk00000001_blk0000006e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011c,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006d
    );
  blk00000001_blk0000006d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011d,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006c
    );
  blk00000001_blk0000006c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011e,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006b
    );
  blk00000001_blk0000006b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000011f,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000006a
    );
  blk00000001_blk0000006a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000120,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000069
    );
  blk00000001_blk00000069 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000121,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000068
    );
  blk00000001_blk00000068 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000122,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000067
    );
  blk00000001_blk00000067 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000123,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000066
    );
  blk00000001_blk00000066 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000124,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000065
    );
  blk00000001_blk00000065 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000125,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000064
    );
  blk00000001_blk00000064 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000126,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000083
    );
  blk00000001_blk00000063 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000127,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000082
    );
  blk00000001_blk00000062 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000128,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000081
    );
  blk00000001_blk00000061 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000129,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000080
    );
  blk00000001_blk00000060 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012a,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007f
    );
  blk00000001_blk0000005f : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012b,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007e
    );
  blk00000001_blk0000005e : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012c,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007d
    );
  blk00000001_blk0000005d : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012d,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007c
    );
  blk00000001_blk0000005c : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012e,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007b
    );
  blk00000001_blk0000005b : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig0000012f,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000007a
    );
  blk00000001_blk0000005a : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000130,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000079
    );
  blk00000001_blk00000059 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000131,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000078
    );
  blk00000001_blk00000058 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000132,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000077
    );
  blk00000001_blk00000057 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000133,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000076
    );
  blk00000001_blk00000056 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000134,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000075
    );
  blk00000001_blk00000055 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig00000112,
      D => blk00000001_sig00000135,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000074
    );
  blk00000001_blk00000021 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(0),
      Q => blk00000001_sig00000105
    );
  blk00000001_blk00000020 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(1),
      Q => blk00000001_sig00000106
    );
  blk00000001_blk0000001f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(2),
      Q => blk00000001_sig00000107
    );
  blk00000001_blk0000001e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(3),
      Q => blk00000001_sig00000108
    );
  blk00000001_blk0000001d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(4),
      Q => blk00000001_sig00000109
    );
  blk00000001_blk0000001c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(5),
      Q => blk00000001_sig0000010a
    );
  blk00000001_blk0000001b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(8),
      Q => blk00000001_sig0000010b
    );
  blk00000001_blk0000001a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(9),
      Q => blk00000001_sig0000010c
    );
  blk00000001_blk00000019 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(10),
      Q => blk00000001_sig0000010d
    );
  blk00000001_blk00000018 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(11),
      Q => blk00000001_sig0000010e
    );
  blk00000001_blk00000017 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(12),
      Q => blk00000001_sig0000010f
    );
  blk00000001_blk00000016 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(13),
      Q => blk00000001_sig00000110
    );
  blk00000001_blk00000015 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => s_axis_config_tdata(14),
      Q => blk00000001_sig00000111
    );
  blk00000001_blk00000014 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000101,
      Q => NlwRenamedSig_OI_s_axis_config_tready
    );
  blk00000001_blk00000013 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig00000102,
      Q => blk00000001_sig00000103
    );
  blk00000001_blk00000012 : FDR
    port map (
      C => aclk,
      D => blk00000001_sig000000da,
      R => blk00000001_sig000000d7,
      Q => blk00000001_sig0000009a
    );
  blk00000001_blk00000011 : FDS
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig000000d7,
      Q => blk00000001_sig000000f7
    );
  blk00000001_blk00000010 : FDS
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000f7,
      S => blk00000001_sig000000d7,
      Q => blk00000001_sig000000f6
    );
  blk00000001_blk0000000f : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000d8,
      R => blk00000001_sig000000f6,
      Q => event_tlast_unexpected
    );
  blk00000001_blk0000000e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000df,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000097
    );
  blk00000001_blk0000000d : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => NlwRenamedSig_OI_m_axis_data_tuser_10_Q,
      S => blk00000001_sig000000f6,
      Q => blk00000001_sig00000099
    );
  blk00000001_blk0000000c : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000db,
      S => blk00000001_sig000000f6,
      Q => blk00000001_sig000000ea
    );
  blk00000001_blk0000000b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig00000096,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000e8
    );
  blk00000001_blk0000000a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000de,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000e7
    );
  blk00000001_blk00000009 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000d9,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000e6
    );
  blk00000001_blk00000008 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000dd,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000e5
    );
  blk00000001_blk00000007 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000dc,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000e9
    );
  blk00000001_blk00000006 : FDR
    port map (
      C => aclk,
      D => blk00000001_sig00000097,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000fa
    );
  blk00000001_blk00000005 : FDRE
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig00000100,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000f3
    );
  blk00000001_blk00000004 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000d3,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000f8
    );
  blk00000001_blk00000003 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_sig000000d2,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig000000f9
    );
  blk00000001_blk00000002 : GND
    port map (
      G => NlwRenamedSig_OI_m_axis_data_tuser_10_Q
    );
  blk00000001_blk00000022_blk00000054 : INV
    port map (
      I => blk00000001_blk00000022_sig000001df,
      O => blk00000001_blk00000022_sig000001f2
    );
  blk00000001_blk00000022_blk00000053 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001df,
      I1 => blk00000001_sig000000f5,
      O => blk00000001_blk00000022_sig00000200
    );
  blk00000001_blk00000022_blk00000052 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001e0,
      I1 => blk00000001_blk00000022_sig000001df,
      I2 => blk00000001_sig000000f5,
      O => blk00000001_blk00000022_sig000001fe
    );
  blk00000001_blk00000022_blk00000051 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001e1,
      I1 => blk00000001_blk00000022_sig000001df,
      I2 => blk00000001_sig000000f5,
      O => blk00000001_blk00000022_sig000001fc
    );
  blk00000001_blk00000022_blk00000050 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001e2,
      I1 => blk00000001_blk00000022_sig000001df,
      I2 => blk00000001_sig000000f5,
      O => blk00000001_blk00000022_sig000001fa
    );
  blk00000001_blk00000022_blk0000004f : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001e3,
      I1 => blk00000001_blk00000022_sig000001df,
      I2 => blk00000001_sig000000f5,
      O => blk00000001_blk00000022_sig000001f8
    );
  blk00000001_blk00000022_blk0000004e : LUT6
    generic map(
      INIT => X"8AAA8A8AAABAAAAA"
    )
    port map (
      I0 => blk00000001_sig00000104,
      I1 => blk00000001_blk00000022_sig00000201,
      I2 => blk00000001_blk00000022_sig000001e0,
      I3 => blk00000001_blk00000022_sig000001df,
      I4 => blk00000001_sig000000f5,
      I5 => blk00000001_sig00000103,
      O => blk00000001_blk00000022_sig000001f1
    );
  blk00000001_blk00000022_blk0000004d : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_blk00000022_sig000001e3,
      I1 => blk00000001_blk00000022_sig000001e1,
      I2 => blk00000001_blk00000022_sig000001e2,
      O => blk00000001_blk00000022_sig00000201
    );
  blk00000001_blk00000022_blk0000004c : XORCY
    port map (
      CI => blk00000001_blk00000022_sig000001ff,
      LI => blk00000001_blk00000022_sig00000200,
      O => blk00000001_blk00000022_sig000001f7
    );
  blk00000001_blk00000022_blk0000004b : XORCY
    port map (
      CI => blk00000001_blk00000022_sig000001fd,
      LI => blk00000001_blk00000022_sig000001fe,
      O => blk00000001_blk00000022_sig000001f6
    );
  blk00000001_blk00000022_blk0000004a : MUXCY
    port map (
      CI => blk00000001_blk00000022_sig000001fd,
      DI => blk00000001_blk00000022_sig000001e0,
      S => blk00000001_blk00000022_sig000001fe,
      O => blk00000001_blk00000022_sig000001ff
    );
  blk00000001_blk00000022_blk00000049 : XORCY
    port map (
      CI => blk00000001_blk00000022_sig000001fb,
      LI => blk00000001_blk00000022_sig000001fc,
      O => blk00000001_blk00000022_sig000001f5
    );
  blk00000001_blk00000022_blk00000048 : MUXCY
    port map (
      CI => blk00000001_blk00000022_sig000001fb,
      DI => blk00000001_blk00000022_sig000001e1,
      S => blk00000001_blk00000022_sig000001fc,
      O => blk00000001_blk00000022_sig000001fd
    );
  blk00000001_blk00000022_blk00000047 : XORCY
    port map (
      CI => blk00000001_blk00000022_sig000001f9,
      LI => blk00000001_blk00000022_sig000001fa,
      O => blk00000001_blk00000022_sig000001f4
    );
  blk00000001_blk00000022_blk00000046 : MUXCY
    port map (
      CI => blk00000001_blk00000022_sig000001f9,
      DI => blk00000001_blk00000022_sig000001e2,
      S => blk00000001_blk00000022_sig000001fa,
      O => blk00000001_blk00000022_sig000001fb
    );
  blk00000001_blk00000022_blk00000045 : XORCY
    port map (
      CI => blk00000001_sig00000103,
      LI => blk00000001_blk00000022_sig000001f8,
      O => blk00000001_blk00000022_sig000001f3
    );
  blk00000001_blk00000022_blk00000044 : MUXCY
    port map (
      CI => blk00000001_sig00000103,
      DI => blk00000001_blk00000022_sig000001e3,
      S => blk00000001_blk00000022_sig000001f8,
      O => blk00000001_blk00000022_sig000001f9
    );
  blk00000001_blk00000022_blk00000043 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000111,
      Q => blk00000001_blk00000022_sig000001e4,
      Q15 => NLW_blk00000001_blk00000022_blk00000043_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000042 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000110,
      Q => blk00000001_blk00000022_sig000001e5,
      Q15 => NLW_blk00000001_blk00000022_blk00000042_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000041 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010f,
      Q => blk00000001_blk00000022_sig000001e6,
      Q15 => NLW_blk00000001_blk00000022_blk00000041_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000040 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010e,
      Q => blk00000001_blk00000022_sig000001e7,
      Q15 => NLW_blk00000001_blk00000022_blk00000040_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010d,
      Q => blk00000001_blk00000022_sig000001e8,
      Q15 => NLW_blk00000001_blk00000022_blk0000003f_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010c,
      Q => blk00000001_blk00000022_sig000001e9,
      Q15 => NLW_blk00000001_blk00000022_blk0000003e_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010b,
      Q => blk00000001_blk00000022_sig000001ea,
      Q15 => NLW_blk00000001_blk00000022_blk0000003d_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig0000010a,
      Q => blk00000001_blk00000022_sig000001eb,
      Q15 => NLW_blk00000001_blk00000022_blk0000003c_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000109,
      Q => blk00000001_blk00000022_sig000001ec,
      Q15 => NLW_blk00000001_blk00000022_blk0000003b_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk0000003a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000108,
      Q => blk00000001_blk00000022_sig000001ed,
      Q15 => NLW_blk00000001_blk00000022_blk0000003a_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000039 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000107,
      Q => blk00000001_blk00000022_sig000001ee,
      Q15 => NLW_blk00000001_blk00000022_blk00000039_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000038 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000106,
      Q => blk00000001_blk00000022_sig000001ef,
      Q15 => NLW_blk00000001_blk00000022_blk00000038_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000037 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000022_sig000001e3,
      A1 => blk00000001_blk00000022_sig000001e2,
      A2 => blk00000001_blk00000022_sig000001e1,
      A3 => blk00000001_blk00000022_sig000001e0,
      CE => blk00000001_sig00000103,
      CLK => aclk,
      D => blk00000001_sig00000105,
      Q => blk00000001_blk00000022_sig000001f0,
      Q15 => NLW_blk00000001_blk00000022_blk00000037_Q15_UNCONNECTED
    );
  blk00000001_blk00000022_blk00000036 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f7,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000022_sig000001df
    );
  blk00000001_blk00000022_blk00000035 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f6,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000022_sig000001e0
    );
  blk00000001_blk00000022_blk00000034 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f5,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000022_sig000001e1
    );
  blk00000001_blk00000022_blk00000033 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f4,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000022_sig000001e2
    );
  blk00000001_blk00000022_blk00000032 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f3,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000022_sig000001e3
    );
  blk00000001_blk00000022_blk00000031 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e4,
      Q => blk00000001_sig00000084
    );
  blk00000001_blk00000022_blk00000030 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e5,
      Q => blk00000001_sig00000085
    );
  blk00000001_blk00000022_blk0000002f : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e6,
      Q => blk00000001_sig00000086
    );
  blk00000001_blk00000022_blk0000002e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e7,
      Q => blk00000001_sig00000087
    );
  blk00000001_blk00000022_blk0000002d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e8,
      Q => blk00000001_sig00000088
    );
  blk00000001_blk00000022_blk0000002c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001e9,
      Q => blk00000001_sig00000089
    );
  blk00000001_blk00000022_blk0000002b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001ea,
      Q => blk00000001_sig00000098
    );
  blk00000001_blk00000022_blk0000002a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001eb,
      Q => blk00000001_sig0000005e
    );
  blk00000001_blk00000022_blk00000029 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001ec,
      Q => blk00000001_sig0000005f
    );
  blk00000001_blk00000022_blk00000028 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001ed,
      Q => blk00000001_sig00000060
    );
  blk00000001_blk00000022_blk00000027 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001ee,
      Q => blk00000001_sig00000061
    );
  blk00000001_blk00000022_blk00000026 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001ef,
      Q => blk00000001_sig00000062
    );
  blk00000001_blk00000022_blk00000025 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f0,
      Q => blk00000001_sig00000063
    );
  blk00000001_blk00000022_blk00000024 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f1,
      S => blk00000001_sig000000f6,
      Q => blk00000001_sig00000104
    );
  blk00000001_blk00000022_blk00000023 : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000022_sig000001f2,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig00000100
    );
  blk00000001_blk000000ba_blk00000116 : INV
    port map (
      I => blk00000001_blk000000ba_sig0000024a,
      O => blk00000001_blk000000ba_sig00000272
    );
  blk00000001_blk000000ba_blk00000115 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024a,
      I1 => blk00000001_sig00000136,
      O => blk00000001_blk000000ba_sig00000280
    );
  blk00000001_blk000000ba_blk00000114 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024b,
      I1 => blk00000001_blk000000ba_sig0000024a,
      I2 => blk00000001_sig00000136,
      O => blk00000001_blk000000ba_sig0000027e
    );
  blk00000001_blk000000ba_blk00000113 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024c,
      I1 => blk00000001_blk000000ba_sig0000024a,
      I2 => blk00000001_sig00000136,
      O => blk00000001_blk000000ba_sig0000027c
    );
  blk00000001_blk000000ba_blk00000112 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024d,
      I1 => blk00000001_blk000000ba_sig0000024a,
      I2 => blk00000001_sig00000136,
      O => blk00000001_blk000000ba_sig0000027a
    );
  blk00000001_blk000000ba_blk00000111 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024e,
      I1 => blk00000001_blk000000ba_sig0000024a,
      I2 => blk00000001_sig00000136,
      O => blk00000001_blk000000ba_sig00000278
    );
  blk00000001_blk000000ba_blk00000110 : LUT6
    generic map(
      INIT => X"8AAA8A8AAABAAAAA"
    )
    port map (
      I0 => blk00000001_sig0000017f,
      I1 => blk00000001_blk000000ba_sig00000282,
      I2 => blk00000001_blk000000ba_sig0000024b,
      I3 => blk00000001_blk000000ba_sig0000024a,
      I4 => blk00000001_sig00000136,
      I5 => blk00000001_sig0000017e,
      O => blk00000001_blk000000ba_sig00000271
    );
  blk00000001_blk000000ba_blk0000010f : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_blk000000ba_sig0000024d,
      I1 => blk00000001_blk000000ba_sig0000024c,
      I2 => blk00000001_blk000000ba_sig0000024e,
      O => blk00000001_blk000000ba_sig00000282
    );
  blk00000001_blk000000ba_blk0000010e : LUT3
    generic map(
      INIT => X"02"
    )
    port map (
      I0 => blk00000001_sig00000136,
      I1 => blk00000001_blk000000ba_sig0000024a,
      I2 => blk00000001_sig000000f6,
      O => blk00000001_blk000000ba_sig00000281
    );
  blk00000001_blk000000ba_blk0000010d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000281,
      Q => blk00000001_sig00000159
    );
  blk00000001_blk000000ba_blk0000010c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig000001a0,
      Q => blk00000001_blk000000ba_sig00000250,
      Q15 => NLW_blk00000001_blk000000ba_blk0000010c_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk0000010b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019f,
      Q => blk00000001_blk000000ba_sig00000251,
      Q15 => NLW_blk00000001_blk000000ba_blk0000010b_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk0000010a : XORCY
    port map (
      CI => blk00000001_blk000000ba_sig0000027f,
      LI => blk00000001_blk000000ba_sig00000280,
      O => blk00000001_blk000000ba_sig00000277
    );
  blk00000001_blk000000ba_blk00000109 : XORCY
    port map (
      CI => blk00000001_blk000000ba_sig0000027d,
      LI => blk00000001_blk000000ba_sig0000027e,
      O => blk00000001_blk000000ba_sig00000276
    );
  blk00000001_blk000000ba_blk00000108 : MUXCY
    port map (
      CI => blk00000001_blk000000ba_sig0000027d,
      DI => blk00000001_blk000000ba_sig0000024b,
      S => blk00000001_blk000000ba_sig0000027e,
      O => blk00000001_blk000000ba_sig0000027f
    );
  blk00000001_blk000000ba_blk00000107 : XORCY
    port map (
      CI => blk00000001_blk000000ba_sig0000027b,
      LI => blk00000001_blk000000ba_sig0000027c,
      O => blk00000001_blk000000ba_sig00000275
    );
  blk00000001_blk000000ba_blk00000106 : MUXCY
    port map (
      CI => blk00000001_blk000000ba_sig0000027b,
      DI => blk00000001_blk000000ba_sig0000024c,
      S => blk00000001_blk000000ba_sig0000027c,
      O => blk00000001_blk000000ba_sig0000027d
    );
  blk00000001_blk000000ba_blk00000105 : XORCY
    port map (
      CI => blk00000001_blk000000ba_sig00000279,
      LI => blk00000001_blk000000ba_sig0000027a,
      O => blk00000001_blk000000ba_sig00000274
    );
  blk00000001_blk000000ba_blk00000104 : MUXCY
    port map (
      CI => blk00000001_blk000000ba_sig00000279,
      DI => blk00000001_blk000000ba_sig0000024d,
      S => blk00000001_blk000000ba_sig0000027a,
      O => blk00000001_blk000000ba_sig0000027b
    );
  blk00000001_blk000000ba_blk00000103 : XORCY
    port map (
      CI => blk00000001_sig0000017e,
      LI => blk00000001_blk000000ba_sig00000278,
      O => blk00000001_blk000000ba_sig00000273
    );
  blk00000001_blk000000ba_blk00000102 : MUXCY
    port map (
      CI => blk00000001_sig0000017e,
      DI => blk00000001_blk000000ba_sig0000024e,
      S => blk00000001_blk000000ba_sig00000278,
      O => blk00000001_blk000000ba_sig00000279
    );
  blk00000001_blk000000ba_blk00000101 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019d,
      Q => blk00000001_blk000000ba_sig00000253,
      Q15 => NLW_blk00000001_blk000000ba_blk00000101_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk00000100 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019c,
      Q => blk00000001_blk000000ba_sig00000254,
      Q15 => NLW_blk00000001_blk000000ba_blk00000100_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ff : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019e,
      Q => blk00000001_blk000000ba_sig00000252,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ff_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000fe : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019a,
      Q => blk00000001_blk000000ba_sig00000256,
      Q15 => NLW_blk00000001_blk000000ba_blk000000fe_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000fd : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000199,
      Q => blk00000001_blk000000ba_sig00000257,
      Q15 => NLW_blk00000001_blk000000ba_blk000000fd_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000fc : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000019b,
      Q => blk00000001_blk000000ba_sig00000255,
      Q15 => NLW_blk00000001_blk000000ba_blk000000fc_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000fb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000198,
      Q => blk00000001_blk000000ba_sig00000258,
      Q15 => NLW_blk00000001_blk000000ba_blk000000fb_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000fa : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000197,
      Q => blk00000001_blk000000ba_sig00000259,
      Q15 => NLW_blk00000001_blk000000ba_blk000000fa_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000196,
      Q => blk00000001_blk000000ba_sig0000025a,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f9_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000195,
      Q => blk00000001_blk000000ba_sig0000025b,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f8_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000193,
      Q => blk00000001_blk000000ba_sig0000025d,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f7_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000192,
      Q => blk00000001_blk000000ba_sig0000025e,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f6_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000194,
      Q => blk00000001_blk000000ba_sig0000025c,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f5_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000190,
      Q => blk00000001_blk000000ba_sig00000260,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f4_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018f,
      Q => blk00000001_blk000000ba_sig00000261,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f3_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f2 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000191,
      Q => blk00000001_blk000000ba_sig0000025f,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f2_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018d,
      Q => blk00000001_blk000000ba_sig00000263,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f1_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000f0 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018c,
      Q => blk00000001_blk000000ba_sig00000264,
      Q15 => NLW_blk00000001_blk000000ba_blk000000f0_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ef : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018e,
      Q => blk00000001_blk000000ba_sig00000262,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ef_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ee : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018b,
      Q => blk00000001_blk000000ba_sig00000265,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ee_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ed : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig0000018a,
      Q => blk00000001_blk000000ba_sig00000266,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ed_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ec : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000189,
      Q => blk00000001_blk000000ba_sig00000267,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ec_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000eb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000188,
      Q => blk00000001_blk000000ba_sig00000268,
      Q15 => NLW_blk00000001_blk000000ba_blk000000eb_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000ea : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000186,
      Q => blk00000001_blk000000ba_sig0000026a,
      Q15 => NLW_blk00000001_blk000000ba_blk000000ea_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000185,
      Q => blk00000001_blk000000ba_sig0000026b,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e9_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e8 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000187,
      Q => blk00000001_blk000000ba_sig00000269,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e8_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000183,
      Q => blk00000001_blk000000ba_sig0000026d,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e7_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e6 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000182,
      Q => blk00000001_blk000000ba_sig0000026e,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e6_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000184,
      Q => blk00000001_blk000000ba_sig0000026c,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e5_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e4 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000180,
      Q => blk00000001_blk000000ba_sig00000270,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e4_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000000ba_sig0000024e,
      A1 => blk00000001_blk000000ba_sig0000024d,
      A2 => blk00000001_blk000000ba_sig0000024c,
      A3 => blk00000001_blk000000ba_sig0000024b,
      CE => blk00000001_sig0000017e,
      CLK => aclk,
      D => blk00000001_sig00000181,
      Q => blk00000001_blk000000ba_sig0000026f,
      Q15 => NLW_blk00000001_blk000000ba_blk000000e3_Q15_UNCONNECTED
    );
  blk00000001_blk000000ba_blk000000e2 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000277,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk000000ba_sig0000024a
    );
  blk00000001_blk000000ba_blk000000e1 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000276,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk000000ba_sig0000024b
    );
  blk00000001_blk000000ba_blk000000e0 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000275,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk000000ba_sig0000024c
    );
  blk00000001_blk000000ba_blk000000df : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000274,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk000000ba_sig0000024d
    );
  blk00000001_blk000000ba_blk000000de : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000273,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk000000ba_sig0000024e
    );
  blk00000001_blk000000ba_blk000000dd : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000250,
      Q => blk00000001_sig0000017b
    );
  blk00000001_blk000000ba_blk000000dc : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000251,
      Q => blk00000001_sig0000017a
    );
  blk00000001_blk000000ba_blk000000db : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000252,
      Q => blk00000001_sig00000179
    );
  blk00000001_blk000000ba_blk000000da : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000253,
      Q => blk00000001_sig00000178
    );
  blk00000001_blk000000ba_blk000000d9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000254,
      Q => blk00000001_sig00000177
    );
  blk00000001_blk000000ba_blk000000d8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000255,
      Q => blk00000001_sig00000176
    );
  blk00000001_blk000000ba_blk000000d7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000256,
      Q => blk00000001_sig00000175
    );
  blk00000001_blk000000ba_blk000000d6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000257,
      Q => blk00000001_sig00000174
    );
  blk00000001_blk000000ba_blk000000d5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000258,
      Q => blk00000001_sig00000173
    );
  blk00000001_blk000000ba_blk000000d4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000259,
      Q => blk00000001_sig00000172
    );
  blk00000001_blk000000ba_blk000000d3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025a,
      Q => blk00000001_sig00000171
    );
  blk00000001_blk000000ba_blk000000d2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025b,
      Q => blk00000001_sig00000170
    );
  blk00000001_blk000000ba_blk000000d1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025c,
      Q => blk00000001_sig0000016f
    );
  blk00000001_blk000000ba_blk000000d0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025d,
      Q => blk00000001_sig0000016e
    );
  blk00000001_blk000000ba_blk000000cf : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025e,
      Q => blk00000001_sig0000016d
    );
  blk00000001_blk000000ba_blk000000ce : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000025f,
      Q => blk00000001_sig0000016c
    );
  blk00000001_blk000000ba_blk000000cd : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000260,
      Q => blk00000001_sig0000016b
    );
  blk00000001_blk000000ba_blk000000cc : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000261,
      Q => blk00000001_sig0000016a
    );
  blk00000001_blk000000ba_blk000000cb : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000262,
      Q => blk00000001_sig00000169
    );
  blk00000001_blk000000ba_blk000000ca : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000263,
      Q => blk00000001_sig00000168
    );
  blk00000001_blk000000ba_blk000000c9 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000264,
      Q => blk00000001_sig00000167
    );
  blk00000001_blk000000ba_blk000000c8 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000265,
      Q => blk00000001_sig00000166
    );
  blk00000001_blk000000ba_blk000000c7 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000266,
      Q => blk00000001_sig00000165
    );
  blk00000001_blk000000ba_blk000000c6 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000267,
      Q => blk00000001_sig00000164
    );
  blk00000001_blk000000ba_blk000000c5 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000268,
      Q => blk00000001_sig00000163
    );
  blk00000001_blk000000ba_blk000000c4 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000269,
      Q => blk00000001_sig00000162
    );
  blk00000001_blk000000ba_blk000000c3 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026a,
      Q => blk00000001_sig00000161
    );
  blk00000001_blk000000ba_blk000000c2 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026b,
      Q => blk00000001_sig00000160
    );
  blk00000001_blk000000ba_blk000000c1 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026c,
      Q => blk00000001_sig0000015f
    );
  blk00000001_blk000000ba_blk000000c0 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026d,
      Q => blk00000001_sig0000015e
    );
  blk00000001_blk000000ba_blk000000bf : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026e,
      Q => blk00000001_sig0000015d
    );
  blk00000001_blk000000ba_blk000000be : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig0000026f,
      Q => blk00000001_sig0000015c
    );
  blk00000001_blk000000ba_blk000000bd : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000270,
      Q => blk00000001_sig0000015b
    );
  blk00000001_blk000000ba_blk000000bc : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000271,
      S => blk00000001_sig000000f6,
      Q => blk00000001_sig0000017f
    );
  blk00000001_blk000000ba_blk000000bb : FDR
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000000ba_sig00000272,
      R => blk00000001_sig000000f6,
      Q => blk00000001_sig0000015a
    );
  blk00000001_blk00000117_blk00000133 : LUT5
    generic map(
      INIT => X"04445544"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      I3 => aclken,
      I4 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig00000292
    );
  blk00000001_blk00000117_blk00000132 : LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      I3 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig00000293
    );
  blk00000001_blk00000117_blk00000131 : LUT6
    generic map(
      INIT => X"4044404440444054"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => blk00000001_sig000000fd,
      I2 => blk00000001_sig000000e1,
      I3 => blk00000001_blk00000117_sig000002a2,
      I4 => blk00000001_blk00000117_sig0000028e,
      I5 => blk00000001_blk00000117_sig000002a4,
      O => blk00000001_blk00000117_sig000002a3
    );
  blk00000001_blk00000117_blk00000130 : LUT3
    generic map(
      INIT => X"7F"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028d,
      I1 => blk00000001_blk00000117_sig0000028c,
      I2 => blk00000001_blk00000117_sig0000028b,
      O => blk00000001_blk00000117_sig000002a4
    );
  blk00000001_blk00000117_blk0000012f : LUT4
    generic map(
      INIT => X"4044"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028a,
      I1 => aclken,
      I2 => m_axis_status_tready,
      I3 => NlwRenamedSig_OI_m_axis_status_tvalid,
      O => blk00000001_blk00000117_sig000002a2
    );
  blk00000001_blk00000117_blk0000012e : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028b,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig00000295
    );
  blk00000001_blk00000117_blk0000012d : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028c,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig00000297
    );
  blk00000001_blk00000117_blk0000012c : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028d,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig00000299
    );
  blk00000001_blk00000117_blk0000012b : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000117_sig0000028e,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I3 => m_axis_status_tready,
      I4 => blk00000001_blk00000117_sig0000028a,
      O => blk00000001_blk00000117_sig0000029b
    );
  blk00000001_blk00000117_blk0000012a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig000002a3,
      Q => blk00000001_sig000000fd
    );
  blk00000001_blk00000117_blk00000129 : LUT3
    generic map(
      INIT => X"A2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_status_tvalid,
      I2 => m_axis_status_tready,
      O => blk00000001_blk00000117_sig00000291
    );
  blk00000001_blk00000117_blk00000128 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000117_sig00000291,
      D => blk00000001_blk00000117_sig000002a1,
      Q => m_axis_status_tdata(0)
    );
  blk00000001_blk00000117_blk00000127 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig000002a0,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000117_sig0000028e
    );
  blk00000001_blk00000117_blk00000126 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig0000029f,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000117_sig0000028d
    );
  blk00000001_blk00000117_blk00000125 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig0000029e,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000117_sig0000028c
    );
  blk00000001_blk00000117_blk00000124 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig0000029d,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000117_sig0000028b
    );
  blk00000001_blk00000117_blk00000123 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig0000029c,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000117_sig0000028a
    );
  blk00000001_blk00000117_blk00000122 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000117_sig0000028e,
      A1 => blk00000001_blk00000117_sig0000028d,
      A2 => blk00000001_blk00000117_sig0000028c,
      A3 => blk00000001_blk00000117_sig0000028b,
      CE => blk00000001_sig000000e1,
      CLK => aclk,
      D => blk00000001_sig000000f4,
      Q => blk00000001_blk00000117_sig000002a1,
      Q15 => NLW_blk00000001_blk00000117_blk00000122_Q15_UNCONNECTED
    );
  blk00000001_blk00000117_blk00000121 : MUXCY
    port map (
      CI => blk00000001_sig000000e1,
      DI => blk00000001_blk00000117_sig0000028e,
      S => blk00000001_blk00000117_sig0000029b,
      O => blk00000001_blk00000117_sig0000029a
    );
  blk00000001_blk00000117_blk00000120 : XORCY
    port map (
      CI => blk00000001_sig000000e1,
      LI => blk00000001_blk00000117_sig0000029b,
      O => blk00000001_blk00000117_sig000002a0
    );
  blk00000001_blk00000117_blk0000011f : MUXCY
    port map (
      CI => blk00000001_blk00000117_sig0000029a,
      DI => blk00000001_blk00000117_sig0000028d,
      S => blk00000001_blk00000117_sig00000299,
      O => blk00000001_blk00000117_sig00000298
    );
  blk00000001_blk00000117_blk0000011e : XORCY
    port map (
      CI => blk00000001_blk00000117_sig0000029a,
      LI => blk00000001_blk00000117_sig00000299,
      O => blk00000001_blk00000117_sig0000029f
    );
  blk00000001_blk00000117_blk0000011d : MUXCY
    port map (
      CI => blk00000001_blk00000117_sig00000298,
      DI => blk00000001_blk00000117_sig0000028c,
      S => blk00000001_blk00000117_sig00000297,
      O => blk00000001_blk00000117_sig00000296
    );
  blk00000001_blk00000117_blk0000011c : XORCY
    port map (
      CI => blk00000001_blk00000117_sig00000298,
      LI => blk00000001_blk00000117_sig00000297,
      O => blk00000001_blk00000117_sig0000029e
    );
  blk00000001_blk00000117_blk0000011b : MUXCY
    port map (
      CI => blk00000001_blk00000117_sig00000296,
      DI => blk00000001_blk00000117_sig0000028b,
      S => blk00000001_blk00000117_sig00000295,
      O => blk00000001_blk00000117_sig00000294
    );
  blk00000001_blk00000117_blk0000011a : XORCY
    port map (
      CI => blk00000001_blk00000117_sig00000296,
      LI => blk00000001_blk00000117_sig00000295,
      O => blk00000001_blk00000117_sig0000029d
    );
  blk00000001_blk00000117_blk00000119 : XORCY
    port map (
      CI => blk00000001_blk00000117_sig00000294,
      LI => blk00000001_blk00000117_sig00000293,
      O => blk00000001_blk00000117_sig0000029c
    );
  blk00000001_blk00000117_blk00000118 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000117_sig00000292,
      Q => NlwRenamedSig_OI_m_axis_status_tvalid
    );
  blk00000001_blk00000134_blk000001a1 : LUT5
    generic map(
      INIT => X"04445544"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      I3 => aclken,
      I4 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig00000303
    );
  blk00000001_blk00000134_blk000001a0 : LUT4
    generic map(
      INIT => X"FFA2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      I3 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig00000304
    );
  blk00000001_blk00000134_blk0000019f : LUT6
    generic map(
      INIT => X"0A0A0A0B000A000A"
    )
    port map (
      I0 => blk00000001_sig000000fc,
      I1 => blk00000001_blk00000134_sig000002fe,
      I2 => blk00000001_sig000000f6,
      I3 => blk00000001_blk00000134_sig0000033b,
      I4 => blk00000001_blk00000134_sig0000033e,
      I5 => blk00000001_sig000000e2,
      O => blk00000001_blk00000134_sig0000033c
    );
  blk00000001_blk00000134_blk0000019e : LUT3
    generic map(
      INIT => X"7F"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fd,
      I1 => blk00000001_blk00000134_sig000002fc,
      I2 => blk00000001_blk00000134_sig000002fb,
      O => blk00000001_blk00000134_sig0000033e
    );
  blk00000001_blk00000134_blk0000019d : LUT4
    generic map(
      INIT => X"4044"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fa,
      I1 => aclken,
      I2 => m_axis_data_tready,
      I3 => NlwRenamedSig_OI_m_axis_data_tvalid,
      O => blk00000001_blk00000134_sig0000033b
    );
  blk00000001_blk00000134_blk0000019c : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fb,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig00000306
    );
  blk00000001_blk00000134_blk0000019b : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fc,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig00000308
    );
  blk00000001_blk00000134_blk0000019a : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fd,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig0000030a
    );
  blk00000001_blk00000134_blk00000199 : LUT5
    generic map(
      INIT => X"AAAA66A6"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fe,
      I1 => aclken,
      I2 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I3 => m_axis_data_tready,
      I4 => blk00000001_blk00000134_sig000002fa,
      O => blk00000001_blk00000134_sig0000030c
    );
  blk00000001_blk00000134_blk00000198 : LUT6
    generic map(
      INIT => X"5455404444444444"
    )
    port map (
      I0 => blk00000001_sig000000f6,
      I1 => blk00000001_sig000000fb,
      I2 => blk00000001_blk00000134_sig000002fa,
      I3 => blk00000001_blk00000134_sig00000302,
      I4 => blk00000001_sig000000e2,
      I5 => blk00000001_blk00000134_sig00000312,
      O => blk00000001_blk00000134_sig0000033d
    );
  blk00000001_blk00000134_blk00000197 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig0000033d,
      Q => blk00000001_sig000000fb
    );
  blk00000001_blk00000134_blk00000196 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig0000033c,
      Q => blk00000001_sig000000fc
    );
  blk00000001_blk00000134_blk00000195 : LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      I0 => blk00000001_blk00000134_sig000002fb,
      I1 => blk00000001_blk00000134_sig000002fc,
      I2 => blk00000001_blk00000134_sig000002fd,
      I3 => blk00000001_blk00000134_sig000002fe,
      O => blk00000001_blk00000134_sig00000312
    );
  blk00000001_blk00000134_blk00000194 : LUT3
    generic map(
      INIT => X"A2"
    )
    port map (
      I0 => aclken,
      I1 => NlwRenamedSig_OI_m_axis_data_tvalid,
      I2 => m_axis_data_tready,
      O => blk00000001_blk00000134_sig00000302
    );
  blk00000001_blk00000134_blk00000193 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000313,
      Q => m_axis_data_tlast
    );
  blk00000001_blk00000134_blk00000192 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000314,
      Q => m_axis_data_tdata(0)
    );
  blk00000001_blk00000134_blk00000191 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000315,
      Q => m_axis_data_tdata(1)
    );
  blk00000001_blk00000134_blk00000190 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000316,
      Q => m_axis_data_tdata(2)
    );
  blk00000001_blk00000134_blk0000018f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000317,
      Q => m_axis_data_tdata(3)
    );
  blk00000001_blk00000134_blk0000018e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000318,
      Q => m_axis_data_tdata(4)
    );
  blk00000001_blk00000134_blk0000018d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000319,
      Q => m_axis_data_tdata(5)
    );
  blk00000001_blk00000134_blk0000018c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031a,
      Q => m_axis_data_tdata(6)
    );
  blk00000001_blk00000134_blk0000018b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031b,
      Q => m_axis_data_tdata(7)
    );
  blk00000001_blk00000134_blk0000018a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031c,
      Q => m_axis_data_tdata(8)
    );
  blk00000001_blk00000134_blk00000189 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031d,
      Q => m_axis_data_tdata(9)
    );
  blk00000001_blk00000134_blk00000188 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031e,
      Q => m_axis_data_tdata(10)
    );
  blk00000001_blk00000134_blk00000187 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000031f,
      Q => m_axis_data_tdata(11)
    );
  blk00000001_blk00000134_blk00000186 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000320,
      Q => m_axis_data_tdata(12)
    );
  blk00000001_blk00000134_blk00000185 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000321,
      Q => m_axis_data_tdata(13)
    );
  blk00000001_blk00000134_blk00000184 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000322,
      Q => m_axis_data_tdata(14)
    );
  blk00000001_blk00000134_blk00000183 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000323,
      Q => m_axis_data_tdata(15)
    );
  blk00000001_blk00000134_blk00000182 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000324,
      Q => m_axis_data_tdata(16)
    );
  blk00000001_blk00000134_blk00000181 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000325,
      Q => m_axis_data_tdata(17)
    );
  blk00000001_blk00000134_blk00000180 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000326,
      Q => m_axis_data_tdata(18)
    );
  blk00000001_blk00000134_blk0000017f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000327,
      Q => m_axis_data_tdata(19)
    );
  blk00000001_blk00000134_blk0000017e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000328,
      Q => m_axis_data_tdata(20)
    );
  blk00000001_blk00000134_blk0000017d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000329,
      Q => m_axis_data_tdata(21)
    );
  blk00000001_blk00000134_blk0000017c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032a,
      Q => m_axis_data_tdata(22)
    );
  blk00000001_blk00000134_blk0000017b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032b,
      Q => m_axis_data_tdata(23)
    );
  blk00000001_blk00000134_blk0000017a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032c,
      Q => m_axis_data_tdata(24)
    );
  blk00000001_blk00000134_blk00000179 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032d,
      Q => m_axis_data_tdata(25)
    );
  blk00000001_blk00000134_blk00000178 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032e,
      Q => m_axis_data_tdata(26)
    );
  blk00000001_blk00000134_blk00000177 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000032f,
      Q => m_axis_data_tdata(27)
    );
  blk00000001_blk00000134_blk00000176 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000330,
      Q => m_axis_data_tdata(28)
    );
  blk00000001_blk00000134_blk00000175 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000331,
      Q => m_axis_data_tdata(29)
    );
  blk00000001_blk00000134_blk00000174 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000332,
      Q => m_axis_data_tdata(30)
    );
  blk00000001_blk00000134_blk00000173 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000333,
      Q => m_axis_data_tdata(31)
    );
  blk00000001_blk00000134_blk00000172 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000334,
      Q => m_axis_data_tuser(0)
    );
  blk00000001_blk00000134_blk00000171 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000335,
      Q => m_axis_data_tuser(1)
    );
  blk00000001_blk00000134_blk00000170 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000336,
      Q => m_axis_data_tuser(2)
    );
  blk00000001_blk00000134_blk0000016f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000337,
      Q => m_axis_data_tuser(3)
    );
  blk00000001_blk00000134_blk0000016e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000338,
      Q => m_axis_data_tuser(4)
    );
  blk00000001_blk00000134_blk0000016d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig00000339,
      Q => m_axis_data_tuser(5)
    );
  blk00000001_blk00000134_blk0000016c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk00000134_sig00000302,
      D => blk00000001_blk00000134_sig0000033a,
      Q => NlwRenamedSig_OI_m_axis_data_tuser_8_Q
    );
  blk00000001_blk00000134_blk0000016b : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig00000311,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000134_sig000002fe
    );
  blk00000001_blk00000134_blk0000016a : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig00000310,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000134_sig000002fd
    );
  blk00000001_blk00000134_blk00000169 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig0000030f,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000134_sig000002fc
    );
  blk00000001_blk00000134_blk00000168 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig0000030e,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000134_sig000002fb
    );
  blk00000001_blk00000134_blk00000167 : FDS
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig0000030d,
      S => blk00000001_sig000000f6,
      Q => blk00000001_blk00000134_sig000002fa
    );
  blk00000001_blk00000134_blk00000166 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000e3,
      Q => blk00000001_blk00000134_sig00000313,
      Q15 => NLW_blk00000001_blk00000134_blk00000166_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000165 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b6,
      Q => blk00000001_blk00000134_sig00000314,
      Q15 => NLW_blk00000001_blk00000134_blk00000165_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000164 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b5,
      Q => blk00000001_blk00000134_sig00000315,
      Q15 => NLW_blk00000001_blk00000134_blk00000164_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000163 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b2,
      Q => blk00000001_blk00000134_sig00000318,
      Q15 => NLW_blk00000001_blk00000134_blk00000163_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000162 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b4,
      Q => blk00000001_blk00000134_sig00000316,
      Q15 => NLW_blk00000001_blk00000134_blk00000162_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000161 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b3,
      Q => blk00000001_blk00000134_sig00000317,
      Q15 => NLW_blk00000001_blk00000134_blk00000161_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000160 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b1,
      Q => blk00000001_blk00000134_sig00000319,
      Q15 => NLW_blk00000001_blk00000134_blk00000160_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b0,
      Q => blk00000001_blk00000134_sig0000031a,
      Q15 => NLW_blk00000001_blk00000134_blk0000015f_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000af,
      Q => blk00000001_blk00000134_sig0000031b,
      Q15 => NLW_blk00000001_blk00000134_blk0000015e_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000ae,
      Q => blk00000001_blk00000134_sig0000031c,
      Q15 => NLW_blk00000001_blk00000134_blk0000015d_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000ab,
      Q => blk00000001_blk00000134_sig0000031f,
      Q15 => NLW_blk00000001_blk00000134_blk0000015c_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000ad,
      Q => blk00000001_blk00000134_sig0000031d,
      Q15 => NLW_blk00000001_blk00000134_blk0000015b_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000015a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000ac,
      Q => blk00000001_blk00000134_sig0000031e,
      Q15 => NLW_blk00000001_blk00000134_blk0000015a_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000159 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000aa,
      Q => blk00000001_blk00000134_sig00000320,
      Q15 => NLW_blk00000001_blk00000134_blk00000159_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000158 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a9,
      Q => blk00000001_blk00000134_sig00000321,
      Q15 => NLW_blk00000001_blk00000134_blk00000158_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000157 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a8,
      Q => blk00000001_blk00000134_sig00000322,
      Q15 => NLW_blk00000001_blk00000134_blk00000157_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000156 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a7,
      Q => blk00000001_blk00000134_sig00000323,
      Q15 => NLW_blk00000001_blk00000134_blk00000156_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000155 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c4,
      Q => blk00000001_blk00000134_sig00000326,
      Q15 => NLW_blk00000001_blk00000134_blk00000155_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000154 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c6,
      Q => blk00000001_blk00000134_sig00000324,
      Q15 => NLW_blk00000001_blk00000134_blk00000154_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000153 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c5,
      Q => blk00000001_blk00000134_sig00000325,
      Q15 => NLW_blk00000001_blk00000134_blk00000153_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000152 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c3,
      Q => blk00000001_blk00000134_sig00000327,
      Q15 => NLW_blk00000001_blk00000134_blk00000152_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000151 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c2,
      Q => blk00000001_blk00000134_sig00000328,
      Q15 => NLW_blk00000001_blk00000134_blk00000151_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000150 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c1,
      Q => blk00000001_blk00000134_sig00000329,
      Q15 => NLW_blk00000001_blk00000134_blk00000150_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000c0,
      Q => blk00000001_blk00000134_sig0000032a,
      Q15 => NLW_blk00000001_blk00000134_blk0000014f_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000bd,
      Q => blk00000001_blk00000134_sig0000032d,
      Q15 => NLW_blk00000001_blk00000134_blk0000014e_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014d : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000bf,
      Q => blk00000001_blk00000134_sig0000032b,
      Q15 => NLW_blk00000001_blk00000134_blk0000014d_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014c : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000be,
      Q => blk00000001_blk00000134_sig0000032c,
      Q15 => NLW_blk00000001_blk00000134_blk0000014c_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000bc,
      Q => blk00000001_blk00000134_sig0000032e,
      Q15 => NLW_blk00000001_blk00000134_blk0000014b_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk0000014a : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000bb,
      Q => blk00000001_blk00000134_sig0000032f,
      Q15 => NLW_blk00000001_blk00000134_blk0000014a_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000149 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000ba,
      Q => blk00000001_blk00000134_sig00000330,
      Q15 => NLW_blk00000001_blk00000134_blk00000149_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000148 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b9,
      Q => blk00000001_blk00000134_sig00000331,
      Q15 => NLW_blk00000001_blk00000134_blk00000148_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000147 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a6,
      Q => blk00000001_blk00000134_sig00000334,
      Q15 => NLW_blk00000001_blk00000134_blk00000147_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000146 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b8,
      Q => blk00000001_blk00000134_sig00000332,
      Q15 => NLW_blk00000001_blk00000134_blk00000146_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000145 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000b7,
      Q => blk00000001_blk00000134_sig00000333,
      Q15 => NLW_blk00000001_blk00000134_blk00000145_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000144 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a5,
      Q => blk00000001_blk00000134_sig00000335,
      Q15 => NLW_blk00000001_blk00000134_blk00000144_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000143 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a4,
      Q => blk00000001_blk00000134_sig00000336,
      Q15 => NLW_blk00000001_blk00000134_blk00000143_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000142 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a3,
      Q => blk00000001_blk00000134_sig00000337,
      Q15 => NLW_blk00000001_blk00000134_blk00000142_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000141 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a2,
      Q => blk00000001_blk00000134_sig00000338,
      Q15 => NLW_blk00000001_blk00000134_blk00000141_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000140 : MUXCY
    port map (
      CI => blk00000001_sig000000e2,
      DI => blk00000001_blk00000134_sig000002fe,
      S => blk00000001_blk00000134_sig0000030c,
      O => blk00000001_blk00000134_sig0000030b
    );
  blk00000001_blk00000134_blk0000013f : XORCY
    port map (
      CI => blk00000001_sig000000e2,
      LI => blk00000001_blk00000134_sig0000030c,
      O => blk00000001_blk00000134_sig00000311
    );
  blk00000001_blk00000134_blk0000013e : MUXCY
    port map (
      CI => blk00000001_blk00000134_sig0000030b,
      DI => blk00000001_blk00000134_sig000002fd,
      S => blk00000001_blk00000134_sig0000030a,
      O => blk00000001_blk00000134_sig00000309
    );
  blk00000001_blk00000134_blk0000013d : XORCY
    port map (
      CI => blk00000001_blk00000134_sig0000030b,
      LI => blk00000001_blk00000134_sig0000030a,
      O => blk00000001_blk00000134_sig00000310
    );
  blk00000001_blk00000134_blk0000013c : MUXCY
    port map (
      CI => blk00000001_blk00000134_sig00000309,
      DI => blk00000001_blk00000134_sig000002fc,
      S => blk00000001_blk00000134_sig00000308,
      O => blk00000001_blk00000134_sig00000307
    );
  blk00000001_blk00000134_blk0000013b : XORCY
    port map (
      CI => blk00000001_blk00000134_sig00000309,
      LI => blk00000001_blk00000134_sig00000308,
      O => blk00000001_blk00000134_sig0000030f
    );
  blk00000001_blk00000134_blk0000013a : MUXCY
    port map (
      CI => blk00000001_blk00000134_sig00000307,
      DI => blk00000001_blk00000134_sig000002fb,
      S => blk00000001_blk00000134_sig00000306,
      O => blk00000001_blk00000134_sig00000305
    );
  blk00000001_blk00000134_blk00000139 : XORCY
    port map (
      CI => blk00000001_blk00000134_sig00000307,
      LI => blk00000001_blk00000134_sig00000306,
      O => blk00000001_blk00000134_sig0000030e
    );
  blk00000001_blk00000134_blk00000138 : XORCY
    port map (
      CI => blk00000001_blk00000134_sig00000305,
      LI => blk00000001_blk00000134_sig00000304,
      O => blk00000001_blk00000134_sig0000030d
    );
  blk00000001_blk00000134_blk00000137 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000a1,
      Q => blk00000001_blk00000134_sig00000339,
      Q15 => NLW_blk00000001_blk00000134_blk00000137_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000136 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk00000134_sig000002fe,
      A1 => blk00000001_blk00000134_sig000002fd,
      A2 => blk00000001_blk00000134_sig000002fc,
      A3 => blk00000001_blk00000134_sig000002fb,
      CE => blk00000001_sig000000e2,
      CLK => aclk,
      D => blk00000001_sig000000cb,
      Q => blk00000001_blk00000134_sig0000033a,
      Q15 => NLW_blk00000001_blk00000134_blk00000136_Q15_UNCONNECTED
    );
  blk00000001_blk00000134_blk00000135 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk00000134_sig00000303,
      Q => NlwRenamedSig_OI_m_axis_data_tvalid
    );
  blk00000001_blk000001a2_blk000001a3_blk00001168 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000efd,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000efd,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000e47,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000e46,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000e45,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000e44,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000e43,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000e42,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000e41,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000e40,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000e3f,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000e3e,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000e3d,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000e3c,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000e3b,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000e3a,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000e39,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000e58,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000e57,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000e56,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000e55,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000e54,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000e53,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000e52,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000e51,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000e50,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000e4f,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000e4e,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000e4d,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000e4c,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000e4b,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000e4a,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000e49,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000efc,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000efb,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000efa,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000ef9,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000ef8,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000ef7,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000ef6,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000ef5,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000ef4,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000ef3,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000ef2,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000ef1,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000ef0,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000eef,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000eee,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000eed,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000eec,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000eeb,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000eea,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000ee9,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000ee8,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000ee7,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000ee6,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000ee5,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000ee4,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000ee3,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000ee2,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000ee1,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000ee0,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000edf,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000ede,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000edd,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000edc,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000edb,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000eda,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000ed9,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000ed8,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000ed7,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000ed6,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000ed5,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000ed4,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000ed3,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000ed2,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000ed1,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000ed0,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000ecf,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000ece,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000ecd,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001168_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001167 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000efc,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000efb,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000efa,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000ef9,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000ef8,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000ef7,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000ef6,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000ef5,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000ef4,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000ef3,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000ef2,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000ef1,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000ef0,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000eef,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000eee,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000eed,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000eec,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000eeb,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000eea,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000ee9,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000ee8,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000ee7,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000ee6,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000ee5,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000ee4,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000ee3,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000ee2,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000ee1,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000ee0,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000edf,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000ede,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000edd,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000edc,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000edb,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000eda,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000ed9,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000ed8,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000ed7,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000ed6,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000ed5,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000ed4,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000ed3,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000ed2,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000ed1,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000ed0,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000ecf,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000ece,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000ecd,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000efe,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000efe,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000e37,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000e36,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000e35,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000e34,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000e33,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000e32,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000e31,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000e30,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000e2f,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000e2e,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000e2d,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000e2c,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000e2b,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000e2a,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000e29,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000c6a,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000c69,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000c68,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000c67,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000c66,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000c65,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000c64,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000c63,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000c62,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000c61,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000c60,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000c5f,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000c5e,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000c5d,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000c5c,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000c5b,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000c5a,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000c59,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000c58,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000c57,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000e69,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000e68,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000e67,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000e66,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000e65,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000e64,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000e63,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000e62,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000e61,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000e60,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000e5f,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000e5e,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000e5d,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000e5c,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000e5b,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000e5a,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001167_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001166 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000e9b,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000e9b,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000dd2,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000dd1,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000dd0,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000dcf,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000dce,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000dcd,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000dcc,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000dcb,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000dca,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000dc9,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000dc8,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000dc7,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000dc6,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000dc5,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000dc4,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000de3,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000de2,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000de1,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000de0,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000ddf,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000dde,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000ddd,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000ddc,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000ddb,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000dda,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000dd9,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000dd8,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000dd7,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000dd6,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000dd5,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000dd4,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000ecc,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000ecb,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000eca,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000ec9,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000ec8,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000ec7,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000ec6,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000ec5,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000ec4,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000ec3,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000ec2,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000ec1,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000ec0,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000ebf,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000ebe,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000ebd,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000ebc,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000ebb,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000eba,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000eb9,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000eb8,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000eb7,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000eb6,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000eb5,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000eb4,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000eb3,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000eb2,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000eb1,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000eb0,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000eaf,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000eae,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000ead,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000eac,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000eab,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000eaa,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000ea9,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000ea8,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000ea7,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000ea6,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000ea5,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000ea4,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000ea3,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000ea2,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000ea1,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000ea0,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000e9f,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000e9e,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000e9d,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001166_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001165 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000ecc,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000ecb,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000eca,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000ec9,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000ec8,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000ec7,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000ec6,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000ec5,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000ec4,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000ec3,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000ec2,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000ec1,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000ec0,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000ebf,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000ebe,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000ebd,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000ebc,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000ebb,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000eba,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000eb9,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000eb8,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000eb7,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000eb6,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000eb5,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000eb4,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000eb3,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000eb2,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000eb1,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000eb0,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000eaf,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000eae,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000ead,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000eac,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000eab,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000eaa,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000ea9,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000ea8,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000ea7,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000ea6,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000ea5,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000ea4,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000ea3,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000ea2,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000ea1,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000ea0,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000e9f,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000e9e,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000e9d,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(0) => blk00000001_blk000001a2_sig00000592,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000dc2,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000dc1,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000dc0,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000dbf,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000dbe,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000dbd,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000dbc,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000dbb,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000dba,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000db9,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000db8,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000db7,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000db6,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000db5,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000db4,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000c92,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000c91,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000c90,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000c8f,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000c8e,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000c8d,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000c8c,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000c8b,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000c8a,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000c89,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000c88,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000c87,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000c86,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000c85,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000c84,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000c83,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000c82,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000c81,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000c80,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000c7f,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000df4,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000df3,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000df2,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000df1,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000df0,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000def,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000dee,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000ded,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000dec,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000deb,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000dea,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000de9,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000de8,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000de7,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000de6,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000de5,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001165_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001164 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000e9b,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000e9b,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000d5f,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000d5e,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000d5d,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000d5c,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000d5b,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000d5a,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000d59,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000d58,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000d57,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000d56,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000d55,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000d54,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000d53,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000d52,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000d51,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000d70,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000d6f,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000d6e,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000d6d,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000d6c,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000d6b,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000d6a,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000d69,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000d68,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000d67,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000d66,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000d65,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000d64,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000d63,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000d62,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000d61,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000e9a,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000e99,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000e98,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000e97,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000e96,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000e95,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000e94,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000e93,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000e92,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000e91,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000e90,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000e8f,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000e8e,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000e8d,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000e8c,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000e8b,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000e8a,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000e89,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000e88,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000e87,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000e86,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000e85,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000e84,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000e83,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000e82,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000e81,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000e80,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000e7f,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000e7e,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000e7d,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000e7c,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000e7b,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000e7a,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000e79,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000e78,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000e77,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000e76,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000e75,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000e74,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000e73,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000e72,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000e71,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000e70,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000e6f,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000e6e,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000e6d,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000e6c,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000e6b,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001164_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001163 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000e9a,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000e99,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000e98,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000e97,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000e96,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000e95,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000e94,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000e93,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000e92,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000e91,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000e90,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000e8f,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000e8e,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000e8d,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000e8c,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000e8b,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000e8a,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000e89,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000e88,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000e87,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000e86,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000e85,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000e84,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000e83,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000e82,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000e81,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000e80,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000e7f,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000e7e,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000e7d,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000e7c,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000e7b,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000e7a,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000e79,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000e78,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000e77,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000e76,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000e75,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000e74,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000e73,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000e72,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000e71,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000e70,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000e6f,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000e6e,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000e6d,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000e6c,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000e6b,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(0) => blk00000001_blk000001a2_sig00000592,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000d4f,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000d4e,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000d4d,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000d4c,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000d4b,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000d4a,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000d49,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000d48,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000d47,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000d46,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000d45,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000d44,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000d43,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000d42,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000d41,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000cba,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000cb9,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000cb8,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000cb7,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000cb6,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000cb5,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000cb4,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000cb3,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000cb2,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000cb1,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000cb0,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000caf,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000cae,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000cad,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000cac,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000cab,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000caa,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000ca9,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000ca8,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000ca7,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000d81,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000d80,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000d7f,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000d7e,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000d7d,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000d7c,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000d7b,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000d7a,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000d79,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000d78,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000d77,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000d76,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000d75,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000d74,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000d73,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000d72,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001163_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001162 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000e28,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000e28,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000e48,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000e47,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000e46,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000e45,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000e44,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000e43,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000e42,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000e41,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000e40,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000e3f,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000e3e,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000e3d,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000e3c,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000e3b,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000e3a,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000e39,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000e6a,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000e69,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000e68,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000e67,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000e66,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000e65,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000e64,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000e63,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000e62,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000e61,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000e60,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000e5f,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000e5e,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000e5d,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000e5c,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000e5b,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000e5a,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000e26,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000e25,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000e24,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000e23,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000e22,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000e21,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000e20,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000e1f,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000e1e,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000e1d,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000e1c,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000e1b,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000e1a,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000e19,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000e18,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000e17,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000e16,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000e15,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000e14,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000e13,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000e12,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000e11,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000e10,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000e0f,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000e0e,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000e0d,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000e0c,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000e0b,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000e0a,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000e09,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000e08,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000e07,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000e06,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000e05,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000e04,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000e03,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000e02,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000e01,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000e00,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000dff,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000dfe,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000dfd,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000dfc,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000dfb,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000dfa,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000df9,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000df8,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000df7,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001162_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001161 : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000e26,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000e25,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000e24,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000e23,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000e22,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000e21,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000e20,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000e1f,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000e1e,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000e1d,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000e1c,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000e1b,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000e1a,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000e19,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000e18,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000e17,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000e16,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000e15,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000e14,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000e13,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000e12,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000e11,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000e10,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000e0f,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000e0e,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000e0d,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000e0c,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000e0b,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000e0a,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000e09,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000e08,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000e07,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000e06,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000e05,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000e04,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000e03,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000e02,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000e01,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000e00,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000dff,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000dfe,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000dfd,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000dfc,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000dfb,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000dfa,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000df9,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000df8,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000df7,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000df6,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000df6,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000e38,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000e37,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000e36,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000e35,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000e34,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000e33,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000e32,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000e31,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000e30,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000e2f,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000e2e,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000e2d,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000e2c,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000e2b,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000e2a,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000e29,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000c7e,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000c7d,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000c7c,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000c7b,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000c7a,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000c79,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000c78,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000c77,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000c76,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000c75,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000c74,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000c73,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000c72,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000c71,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000c70,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000c6f,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000c6e,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000c6d,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000c6c,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000c6b,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000e59,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000e58,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000e57,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000e56,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000e55,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000e54,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000e53,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000e52,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000e51,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000e50,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000e4f,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000e4e,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000e4d,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000e4c,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000e4b,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000e4a,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000e49,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001161_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001160 : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(0) => blk00000001_blk000001a2_sig00000592,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000dd3,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000dd2,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000dd1,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000dd0,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000dcf,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000dce,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000dcd,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000dcc,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000dcb,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000dca,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000dc9,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000dc8,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000dc7,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000dc6,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000dc5,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000dc4,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000df5,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000df4,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000df3,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000df2,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000df1,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000df0,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000def,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000dee,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000ded,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000dec,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000deb,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000dea,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000de9,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000de8,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000de7,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000de6,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000de5,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000db3,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000db2,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000db1,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000db0,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000daf,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000dae,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000dad,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000dac,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000dab,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000daa,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000da9,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000da8,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000da7,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000da6,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000da5,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000da4,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000da3,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000da2,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000da1,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000da0,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000d9f,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000d9e,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000d9d,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000d9c,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000d9b,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000d9a,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000d99,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000d98,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000d97,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000d96,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000d95,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000d94,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000d93,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000d92,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000d91,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000d90,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000d8f,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000d8e,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000d8d,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000d8c,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000d8b,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000d8a,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000d89,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000d88,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000d87,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000d86,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000d85,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000d84,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001160_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115f : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000db3,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000db2,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000db1,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000db0,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000daf,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000dae,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000dad,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000dac,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000dab,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000daa,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000da9,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000da8,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000da7,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000da6,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000da5,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000da4,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000da3,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000da2,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000da1,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000da0,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000d9f,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000d9e,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000d9d,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000d9c,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000d9b,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000d9a,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000d99,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000d98,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000d97,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000d96,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000d95,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000d94,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000d93,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000d92,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000d91,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000d90,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000d8f,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000d8e,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000d8d,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000d8c,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000d8b,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000d8a,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000d89,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000d88,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000d87,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000d86,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000d85,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000d84,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000d83,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000d83,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000dc3,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000dc2,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000dc1,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000dc0,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000dbf,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000dbe,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000dbd,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000dbc,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000dbb,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000dba,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000db9,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000db8,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000db7,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000db6,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000db5,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000db4,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000ca6,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000ca5,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000ca4,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000ca3,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000ca2,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000ca1,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000ca0,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000c9f,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000c9e,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000c9d,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000c9c,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000c9b,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000c9a,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000c99,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000c98,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000c97,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000c96,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000c95,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000c94,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000c93,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000de4,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000de3,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000de2,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000de1,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000de0,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000ddf,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000dde,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000ddd,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000ddc,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000ddb,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000dda,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000dd9,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000dd8,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000dd7,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000dd6,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000dd5,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000dd4,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115f_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115e : DSP48E
    generic map(
      ACASCREG => 1,
      ALUMODEREG => 1,
      AREG => 1,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 1,
      BREG => 1,
      B_INPUT => "DIRECT",
      CARRYINREG => 1,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_blk000001a2_sig00000592,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_blk000001a2_sig00000592,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(0) => blk00000001_blk000001a2_sig00000592,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000d60,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000d5f,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000d5e,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000d5d,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000d5c,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000d5b,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000d5a,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000d59,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000d58,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000d57,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000d56,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000d55,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000d54,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000d53,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000d52,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000d51,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000d82,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000d81,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000d80,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000d7f,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000d7e,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000d7d,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000d7c,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000d7b,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000d7a,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000d79,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000d78,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000d77,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000d76,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000d75,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000d74,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000d73,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000d72,
      PCOUT(47) => blk00000001_blk000001a2_blk000001a3_sig00000d3f,
      PCOUT(46) => blk00000001_blk000001a2_blk000001a3_sig00000d3e,
      PCOUT(45) => blk00000001_blk000001a2_blk000001a3_sig00000d3d,
      PCOUT(44) => blk00000001_blk000001a2_blk000001a3_sig00000d3c,
      PCOUT(43) => blk00000001_blk000001a2_blk000001a3_sig00000d3b,
      PCOUT(42) => blk00000001_blk000001a2_blk000001a3_sig00000d3a,
      PCOUT(41) => blk00000001_blk000001a2_blk000001a3_sig00000d39,
      PCOUT(40) => blk00000001_blk000001a2_blk000001a3_sig00000d38,
      PCOUT(39) => blk00000001_blk000001a2_blk000001a3_sig00000d37,
      PCOUT(38) => blk00000001_blk000001a2_blk000001a3_sig00000d36,
      PCOUT(37) => blk00000001_blk000001a2_blk000001a3_sig00000d35,
      PCOUT(36) => blk00000001_blk000001a2_blk000001a3_sig00000d34,
      PCOUT(35) => blk00000001_blk000001a2_blk000001a3_sig00000d33,
      PCOUT(34) => blk00000001_blk000001a2_blk000001a3_sig00000d32,
      PCOUT(33) => blk00000001_blk000001a2_blk000001a3_sig00000d31,
      PCOUT(32) => blk00000001_blk000001a2_blk000001a3_sig00000d30,
      PCOUT(31) => blk00000001_blk000001a2_blk000001a3_sig00000d2f,
      PCOUT(30) => blk00000001_blk000001a2_blk000001a3_sig00000d2e,
      PCOUT(29) => blk00000001_blk000001a2_blk000001a3_sig00000d2d,
      PCOUT(28) => blk00000001_blk000001a2_blk000001a3_sig00000d2c,
      PCOUT(27) => blk00000001_blk000001a2_blk000001a3_sig00000d2b,
      PCOUT(26) => blk00000001_blk000001a2_blk000001a3_sig00000d2a,
      PCOUT(25) => blk00000001_blk000001a2_blk000001a3_sig00000d29,
      PCOUT(24) => blk00000001_blk000001a2_blk000001a3_sig00000d28,
      PCOUT(23) => blk00000001_blk000001a2_blk000001a3_sig00000d27,
      PCOUT(22) => blk00000001_blk000001a2_blk000001a3_sig00000d26,
      PCOUT(21) => blk00000001_blk000001a2_blk000001a3_sig00000d25,
      PCOUT(20) => blk00000001_blk000001a2_blk000001a3_sig00000d24,
      PCOUT(19) => blk00000001_blk000001a2_blk000001a3_sig00000d23,
      PCOUT(18) => blk00000001_blk000001a2_blk000001a3_sig00000d22,
      PCOUT(17) => blk00000001_blk000001a2_blk000001a3_sig00000d21,
      PCOUT(16) => blk00000001_blk000001a2_blk000001a3_sig00000d20,
      PCOUT(15) => blk00000001_blk000001a2_blk000001a3_sig00000d1f,
      PCOUT(14) => blk00000001_blk000001a2_blk000001a3_sig00000d1e,
      PCOUT(13) => blk00000001_blk000001a2_blk000001a3_sig00000d1d,
      PCOUT(12) => blk00000001_blk000001a2_blk000001a3_sig00000d1c,
      PCOUT(11) => blk00000001_blk000001a2_blk000001a3_sig00000d1b,
      PCOUT(10) => blk00000001_blk000001a2_blk000001a3_sig00000d1a,
      PCOUT(9) => blk00000001_blk000001a2_blk000001a3_sig00000d19,
      PCOUT(8) => blk00000001_blk000001a2_blk000001a3_sig00000d18,
      PCOUT(7) => blk00000001_blk000001a2_blk000001a3_sig00000d17,
      PCOUT(6) => blk00000001_blk000001a2_blk000001a3_sig00000d16,
      PCOUT(5) => blk00000001_blk000001a2_blk000001a3_sig00000d15,
      PCOUT(4) => blk00000001_blk000001a2_blk000001a3_sig00000d14,
      PCOUT(3) => blk00000001_blk000001a2_blk000001a3_sig00000d13,
      PCOUT(2) => blk00000001_blk000001a2_blk000001a3_sig00000d12,
      PCOUT(1) => blk00000001_blk000001a2_blk000001a3_sig00000d11,
      PCOUT(0) => blk00000001_blk000001a2_blk000001a3_sig00000d10,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_sig00000592,
      PCIN(46) => blk00000001_blk000001a2_sig00000592,
      PCIN(45) => blk00000001_blk000001a2_sig00000592,
      PCIN(44) => blk00000001_blk000001a2_sig00000592,
      PCIN(43) => blk00000001_blk000001a2_sig00000592,
      PCIN(42) => blk00000001_blk000001a2_sig00000592,
      PCIN(41) => blk00000001_blk000001a2_sig00000592,
      PCIN(40) => blk00000001_blk000001a2_sig00000592,
      PCIN(39) => blk00000001_blk000001a2_sig00000592,
      PCIN(38) => blk00000001_blk000001a2_sig00000592,
      PCIN(37) => blk00000001_blk000001a2_sig00000592,
      PCIN(36) => blk00000001_blk000001a2_sig00000592,
      PCIN(35) => blk00000001_blk000001a2_sig00000592,
      PCIN(34) => blk00000001_blk000001a2_sig00000592,
      PCIN(33) => blk00000001_blk000001a2_sig00000592,
      PCIN(32) => blk00000001_blk000001a2_sig00000592,
      PCIN(31) => blk00000001_blk000001a2_sig00000592,
      PCIN(30) => blk00000001_blk000001a2_sig00000592,
      PCIN(29) => blk00000001_blk000001a2_sig00000592,
      PCIN(28) => blk00000001_blk000001a2_sig00000592,
      PCIN(27) => blk00000001_blk000001a2_sig00000592,
      PCIN(26) => blk00000001_blk000001a2_sig00000592,
      PCIN(25) => blk00000001_blk000001a2_sig00000592,
      PCIN(24) => blk00000001_blk000001a2_sig00000592,
      PCIN(23) => blk00000001_blk000001a2_sig00000592,
      PCIN(22) => blk00000001_blk000001a2_sig00000592,
      PCIN(21) => blk00000001_blk000001a2_sig00000592,
      PCIN(20) => blk00000001_blk000001a2_sig00000592,
      PCIN(19) => blk00000001_blk000001a2_sig00000592,
      PCIN(18) => blk00000001_blk000001a2_sig00000592,
      PCIN(17) => blk00000001_blk000001a2_sig00000592,
      PCIN(16) => blk00000001_blk000001a2_sig00000592,
      PCIN(15) => blk00000001_blk000001a2_sig00000592,
      PCIN(14) => blk00000001_blk000001a2_sig00000592,
      PCIN(13) => blk00000001_blk000001a2_sig00000592,
      PCIN(12) => blk00000001_blk000001a2_sig00000592,
      PCIN(11) => blk00000001_blk000001a2_sig00000592,
      PCIN(10) => blk00000001_blk000001a2_sig00000592,
      PCIN(9) => blk00000001_blk000001a2_sig00000592,
      PCIN(8) => blk00000001_blk000001a2_sig00000592,
      PCIN(7) => blk00000001_blk000001a2_sig00000592,
      PCIN(6) => blk00000001_blk000001a2_sig00000592,
      PCIN(5) => blk00000001_blk000001a2_sig00000592,
      PCIN(4) => blk00000001_blk000001a2_sig00000592,
      PCIN(3) => blk00000001_blk000001a2_sig00000592,
      PCIN(2) => blk00000001_blk000001a2_sig00000592,
      PCIN(1) => blk00000001_blk000001a2_sig00000592,
      PCIN(0) => blk00000001_blk000001a2_sig00000592,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_BCOUT_0_UNCONNECTED,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_32_UNCONNECTED,
      P(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_31_UNCONNECTED,
      P(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_30_UNCONNECTED,
      P(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_29_UNCONNECTED,
      P(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_28_UNCONNECTED,
      P(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_27_UNCONNECTED,
      P(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_26_UNCONNECTED,
      P(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_25_UNCONNECTED,
      P(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_24_UNCONNECTED,
      P(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_23_UNCONNECTED,
      P(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_22_UNCONNECTED,
      P(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_21_UNCONNECTED,
      P(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_20_UNCONNECTED,
      P(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_19_UNCONNECTED,
      P(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_18_UNCONNECTED,
      P(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_17_UNCONNECTED,
      P(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_16_UNCONNECTED,
      P(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_15_UNCONNECTED,
      P(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_14_UNCONNECTED,
      P(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_13_UNCONNECTED,
      P(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_12_UNCONNECTED,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115e_P_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115d : DSP48E
    generic map(
      ACASCREG => 2,
      ALUMODEREG => 1,
      AREG => 2,
      AUTORESET_PATTERN_DETECT => FALSE,
      AUTORESET_PATTERN_DETECT_OPTINV => "MATCH",
      A_INPUT => "DIRECT",
      BCASCREG => 2,
      BREG => 2,
      B_INPUT => "DIRECT",
      CARRYINREG => 0,
      CARRYINSELREG => 0,
      CREG => 0,
      MASK => X"000000000000",
      MREG => 1,
      MULTCARRYINREG => 0,
      OPMODEREG => 0,
      PATTERN => X"000000000000",
      PREG => 1,
      SEL_MASK => "MASK",
      SEL_PATTERN => "PATTERN",
      SEL_ROUNDING_MASK => "SEL_MASK",
      SIM_MODE => "SAFE",
      USE_MULT => "MULT_S",
      USE_PATTERN_DETECT => "NO_PATDET",
      USE_SIMD => "ONE48"
    )
    port map (
      CEM => blk00000001_sig0000009a,
      CLK => aclk,
      PATTERNBDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PATTERNBDETECT_UNCONNECTED,
      RSTC => blk00000001_blk000001a2_sig00000592,
      CEB1 => blk00000001_sig0000009a,
      MULTSIGNOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_MULTSIGNOUT_UNCONNECTED,
      CEC => blk00000001_blk000001a2_sig00000592,
      RSTM => blk00000001_blk000001a2_sig00000592,
      MULTSIGNIN => blk00000001_blk000001a2_sig00000592,
      CEB2 => blk00000001_sig0000009a,
      RSTCTRL => blk00000001_blk000001a2_sig00000592,
      CEP => blk00000001_sig0000009a,
      CARRYCASCOUT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYCASCOUT_UNCONNECTED,
      RSTA => blk00000001_blk000001a2_sig00000592,
      CECARRYIN => blk00000001_blk000001a2_sig00000592,
      UNDERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_UNDERFLOW_UNCONNECTED,
      PATTERNDETECT => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PATTERNDETECT_UNCONNECTED,
      RSTALUMODE => blk00000001_blk000001a2_sig00000592,
      RSTALLCARRYIN => blk00000001_blk000001a2_sig00000592,
      CEALUMODE => blk00000001_sig0000009a,
      CEA2 => blk00000001_sig0000009a,
      CEA1 => blk00000001_sig0000009a,
      RSTB => blk00000001_blk000001a2_sig00000592,
      CEMULTCARRYIN => blk00000001_blk000001a2_sig00000592,
      OVERFLOW => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_OVERFLOW_UNCONNECTED,
      CECTRL => blk00000001_blk000001a2_sig00000592,
      CARRYIN => blk00000001_blk000001a2_sig00000592,
      CARRYCASCIN => blk00000001_blk000001a2_sig00000592,
      RSTP => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(2) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(1) => blk00000001_blk000001a2_sig00000592,
      CARRYINSEL(0) => blk00000001_blk000001a2_sig00000592,
      C(47) => blk00000001_blk000001a2_sig00000592,
      C(46) => blk00000001_blk000001a2_sig00000592,
      C(45) => blk00000001_blk000001a2_sig00000592,
      C(44) => blk00000001_blk000001a2_sig00000592,
      C(43) => blk00000001_blk000001a2_sig00000592,
      C(42) => blk00000001_blk000001a2_sig00000592,
      C(41) => blk00000001_blk000001a2_sig00000592,
      C(40) => blk00000001_blk000001a2_sig00000592,
      C(39) => blk00000001_blk000001a2_sig00000592,
      C(38) => blk00000001_blk000001a2_sig00000592,
      C(37) => blk00000001_blk000001a2_sig00000592,
      C(36) => blk00000001_blk000001a2_sig00000592,
      C(35) => blk00000001_blk000001a2_sig00000592,
      C(34) => blk00000001_blk000001a2_sig00000592,
      C(33) => blk00000001_blk000001a2_sig00000592,
      C(32) => blk00000001_blk000001a2_sig00000592,
      C(31) => blk00000001_blk000001a2_sig00000592,
      C(30) => blk00000001_blk000001a2_sig00000592,
      C(29) => blk00000001_blk000001a2_sig00000592,
      C(28) => blk00000001_blk000001a2_sig00000592,
      C(27) => blk00000001_blk000001a2_sig00000592,
      C(26) => blk00000001_blk000001a2_sig00000592,
      C(25) => blk00000001_blk000001a2_sig00000592,
      C(24) => blk00000001_blk000001a2_sig00000592,
      C(23) => blk00000001_blk000001a2_sig00000592,
      C(22) => blk00000001_blk000001a2_sig00000592,
      C(21) => blk00000001_blk000001a2_sig00000592,
      C(20) => blk00000001_blk000001a2_sig00000592,
      C(19) => blk00000001_blk000001a2_sig00000592,
      C(18) => blk00000001_blk000001a2_sig00000592,
      C(17) => blk00000001_blk000001a2_sig00000592,
      C(16) => blk00000001_blk000001a2_sig00000592,
      C(15) => blk00000001_blk000001a2_sig00000592,
      C(14) => blk00000001_blk000001a2_sig00000592,
      C(13) => blk00000001_blk000001a2_sig00000592,
      C(12) => blk00000001_blk000001a2_sig00000592,
      C(11) => blk00000001_blk000001a2_sig00000592,
      C(10) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(8) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(7) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(6) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(5) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      C(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      PCIN(47) => blk00000001_blk000001a2_blk000001a3_sig00000d3f,
      PCIN(46) => blk00000001_blk000001a2_blk000001a3_sig00000d3e,
      PCIN(45) => blk00000001_blk000001a2_blk000001a3_sig00000d3d,
      PCIN(44) => blk00000001_blk000001a2_blk000001a3_sig00000d3c,
      PCIN(43) => blk00000001_blk000001a2_blk000001a3_sig00000d3b,
      PCIN(42) => blk00000001_blk000001a2_blk000001a3_sig00000d3a,
      PCIN(41) => blk00000001_blk000001a2_blk000001a3_sig00000d39,
      PCIN(40) => blk00000001_blk000001a2_blk000001a3_sig00000d38,
      PCIN(39) => blk00000001_blk000001a2_blk000001a3_sig00000d37,
      PCIN(38) => blk00000001_blk000001a2_blk000001a3_sig00000d36,
      PCIN(37) => blk00000001_blk000001a2_blk000001a3_sig00000d35,
      PCIN(36) => blk00000001_blk000001a2_blk000001a3_sig00000d34,
      PCIN(35) => blk00000001_blk000001a2_blk000001a3_sig00000d33,
      PCIN(34) => blk00000001_blk000001a2_blk000001a3_sig00000d32,
      PCIN(33) => blk00000001_blk000001a2_blk000001a3_sig00000d31,
      PCIN(32) => blk00000001_blk000001a2_blk000001a3_sig00000d30,
      PCIN(31) => blk00000001_blk000001a2_blk000001a3_sig00000d2f,
      PCIN(30) => blk00000001_blk000001a2_blk000001a3_sig00000d2e,
      PCIN(29) => blk00000001_blk000001a2_blk000001a3_sig00000d2d,
      PCIN(28) => blk00000001_blk000001a2_blk000001a3_sig00000d2c,
      PCIN(27) => blk00000001_blk000001a2_blk000001a3_sig00000d2b,
      PCIN(26) => blk00000001_blk000001a2_blk000001a3_sig00000d2a,
      PCIN(25) => blk00000001_blk000001a2_blk000001a3_sig00000d29,
      PCIN(24) => blk00000001_blk000001a2_blk000001a3_sig00000d28,
      PCIN(23) => blk00000001_blk000001a2_blk000001a3_sig00000d27,
      PCIN(22) => blk00000001_blk000001a2_blk000001a3_sig00000d26,
      PCIN(21) => blk00000001_blk000001a2_blk000001a3_sig00000d25,
      PCIN(20) => blk00000001_blk000001a2_blk000001a3_sig00000d24,
      PCIN(19) => blk00000001_blk000001a2_blk000001a3_sig00000d23,
      PCIN(18) => blk00000001_blk000001a2_blk000001a3_sig00000d22,
      PCIN(17) => blk00000001_blk000001a2_blk000001a3_sig00000d21,
      PCIN(16) => blk00000001_blk000001a2_blk000001a3_sig00000d20,
      PCIN(15) => blk00000001_blk000001a2_blk000001a3_sig00000d1f,
      PCIN(14) => blk00000001_blk000001a2_blk000001a3_sig00000d1e,
      PCIN(13) => blk00000001_blk000001a2_blk000001a3_sig00000d1d,
      PCIN(12) => blk00000001_blk000001a2_blk000001a3_sig00000d1c,
      PCIN(11) => blk00000001_blk000001a2_blk000001a3_sig00000d1b,
      PCIN(10) => blk00000001_blk000001a2_blk000001a3_sig00000d1a,
      PCIN(9) => blk00000001_blk000001a2_blk000001a3_sig00000d19,
      PCIN(8) => blk00000001_blk000001a2_blk000001a3_sig00000d18,
      PCIN(7) => blk00000001_blk000001a2_blk000001a3_sig00000d17,
      PCIN(6) => blk00000001_blk000001a2_blk000001a3_sig00000d16,
      PCIN(5) => blk00000001_blk000001a2_blk000001a3_sig00000d15,
      PCIN(4) => blk00000001_blk000001a2_blk000001a3_sig00000d14,
      PCIN(3) => blk00000001_blk000001a2_blk000001a3_sig00000d13,
      PCIN(2) => blk00000001_blk000001a2_blk000001a3_sig00000d12,
      PCIN(1) => blk00000001_blk000001a2_blk000001a3_sig00000d11,
      PCIN(0) => blk00000001_blk000001a2_blk000001a3_sig00000d10,
      ALUMODE(3) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(2) => blk00000001_blk000001a2_sig00000592,
      ALUMODE(1) => blk00000001_blk000001a2_blk000001a3_sig00000d0f,
      ALUMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000d0f,
      B(17) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(16) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(15) => blk00000001_blk000001a2_blk000001a3_sig00000d50,
      B(14) => blk00000001_blk000001a2_blk000001a3_sig00000d4f,
      B(13) => blk00000001_blk000001a2_blk000001a3_sig00000d4e,
      B(12) => blk00000001_blk000001a2_blk000001a3_sig00000d4d,
      B(11) => blk00000001_blk000001a2_blk000001a3_sig00000d4c,
      B(10) => blk00000001_blk000001a2_blk000001a3_sig00000d4b,
      B(9) => blk00000001_blk000001a2_blk000001a3_sig00000d4a,
      B(8) => blk00000001_blk000001a2_blk000001a3_sig00000d49,
      B(7) => blk00000001_blk000001a2_blk000001a3_sig00000d48,
      B(6) => blk00000001_blk000001a2_blk000001a3_sig00000d47,
      B(5) => blk00000001_blk000001a2_blk000001a3_sig00000d46,
      B(4) => blk00000001_blk000001a2_blk000001a3_sig00000d45,
      B(3) => blk00000001_blk000001a2_blk000001a3_sig00000d44,
      B(2) => blk00000001_blk000001a2_blk000001a3_sig00000d43,
      B(1) => blk00000001_blk000001a2_blk000001a3_sig00000d42,
      B(0) => blk00000001_blk000001a2_blk000001a3_sig00000d41,
      P(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_47_UNCONNECTED,
      P(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_46_UNCONNECTED,
      P(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_45_UNCONNECTED,
      P(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_44_UNCONNECTED,
      P(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_43_UNCONNECTED,
      P(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_42_UNCONNECTED,
      P(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_41_UNCONNECTED,
      P(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_40_UNCONNECTED,
      P(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_39_UNCONNECTED,
      P(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_38_UNCONNECTED,
      P(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_37_UNCONNECTED,
      P(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_36_UNCONNECTED,
      P(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_35_UNCONNECTED,
      P(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_34_UNCONNECTED,
      P(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_33_UNCONNECTED,
      P(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_32_UNCONNECTED,
      P(31) => blk00000001_blk000001a2_blk000001a3_sig00000cce,
      P(30) => blk00000001_blk000001a2_blk000001a3_sig00000ccd,
      P(29) => blk00000001_blk000001a2_blk000001a3_sig00000ccc,
      P(28) => blk00000001_blk000001a2_blk000001a3_sig00000ccb,
      P(27) => blk00000001_blk000001a2_blk000001a3_sig00000cca,
      P(26) => blk00000001_blk000001a2_blk000001a3_sig00000cc9,
      P(25) => blk00000001_blk000001a2_blk000001a3_sig00000cc8,
      P(24) => blk00000001_blk000001a2_blk000001a3_sig00000cc7,
      P(23) => blk00000001_blk000001a2_blk000001a3_sig00000cc6,
      P(22) => blk00000001_blk000001a2_blk000001a3_sig00000cc5,
      P(21) => blk00000001_blk000001a2_blk000001a3_sig00000cc4,
      P(20) => blk00000001_blk000001a2_blk000001a3_sig00000cc3,
      P(19) => blk00000001_blk000001a2_blk000001a3_sig00000cc2,
      P(18) => blk00000001_blk000001a2_blk000001a3_sig00000cc1,
      P(17) => blk00000001_blk000001a2_blk000001a3_sig00000cc0,
      P(16) => blk00000001_blk000001a2_blk000001a3_sig00000cbf,
      P(15) => blk00000001_blk000001a2_blk000001a3_sig00000cbe,
      P(14) => blk00000001_blk000001a2_blk000001a3_sig00000cbd,
      P(13) => blk00000001_blk000001a2_blk000001a3_sig00000cbc,
      P(12) => blk00000001_blk000001a2_blk000001a3_sig00000cbb,
      P(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_11_UNCONNECTED,
      P(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_10_UNCONNECTED,
      P(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_9_UNCONNECTED,
      P(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_8_UNCONNECTED,
      P(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_7_UNCONNECTED,
      P(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_6_UNCONNECTED,
      P(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_5_UNCONNECTED,
      P(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_4_UNCONNECTED,
      P(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_3_UNCONNECTED,
      P(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_2_UNCONNECTED,
      P(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_1_UNCONNECTED,
      P(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_P_0_UNCONNECTED,
      A(29) => blk00000001_blk000001a2_sig00000592,
      A(28) => blk00000001_blk000001a2_sig00000592,
      A(27) => blk00000001_blk000001a2_sig00000592,
      A(26) => blk00000001_blk000001a2_sig00000592,
      A(25) => blk00000001_blk000001a2_sig00000592,
      A(24) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(23) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(22) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(21) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(20) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(19) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(18) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(17) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(16) => blk00000001_blk000001a2_blk000001a3_sig00000d71,
      A(15) => blk00000001_blk000001a2_blk000001a3_sig00000d70,
      A(14) => blk00000001_blk000001a2_blk000001a3_sig00000d6f,
      A(13) => blk00000001_blk000001a2_blk000001a3_sig00000d6e,
      A(12) => blk00000001_blk000001a2_blk000001a3_sig00000d6d,
      A(11) => blk00000001_blk000001a2_blk000001a3_sig00000d6c,
      A(10) => blk00000001_blk000001a2_blk000001a3_sig00000d6b,
      A(9) => blk00000001_blk000001a2_blk000001a3_sig00000d6a,
      A(8) => blk00000001_blk000001a2_blk000001a3_sig00000d69,
      A(7) => blk00000001_blk000001a2_blk000001a3_sig00000d68,
      A(6) => blk00000001_blk000001a2_blk000001a3_sig00000d67,
      A(5) => blk00000001_blk000001a2_blk000001a3_sig00000d66,
      A(4) => blk00000001_blk000001a2_blk000001a3_sig00000d65,
      A(3) => blk00000001_blk000001a2_blk000001a3_sig00000d64,
      A(2) => blk00000001_blk000001a2_blk000001a3_sig00000d63,
      A(1) => blk00000001_blk000001a2_blk000001a3_sig00000d62,
      A(0) => blk00000001_blk000001a2_blk000001a3_sig00000d61,
      PCOUT(47) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_47_UNCONNECTED,
      PCOUT(46) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_46_UNCONNECTED,
      PCOUT(45) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_45_UNCONNECTED,
      PCOUT(44) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_44_UNCONNECTED,
      PCOUT(43) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_43_UNCONNECTED,
      PCOUT(42) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_42_UNCONNECTED,
      PCOUT(41) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_41_UNCONNECTED,
      PCOUT(40) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_40_UNCONNECTED,
      PCOUT(39) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_39_UNCONNECTED,
      PCOUT(38) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_38_UNCONNECTED,
      PCOUT(37) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_37_UNCONNECTED,
      PCOUT(36) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_36_UNCONNECTED,
      PCOUT(35) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_35_UNCONNECTED,
      PCOUT(34) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_34_UNCONNECTED,
      PCOUT(33) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_33_UNCONNECTED,
      PCOUT(32) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_32_UNCONNECTED,
      PCOUT(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_31_UNCONNECTED,
      PCOUT(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_30_UNCONNECTED,
      PCOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_29_UNCONNECTED,
      PCOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_28_UNCONNECTED,
      PCOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_27_UNCONNECTED,
      PCOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_26_UNCONNECTED,
      PCOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_25_UNCONNECTED,
      PCOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_24_UNCONNECTED,
      PCOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_23_UNCONNECTED,
      PCOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_22_UNCONNECTED,
      PCOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_21_UNCONNECTED,
      PCOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_20_UNCONNECTED,
      PCOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_19_UNCONNECTED,
      PCOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_18_UNCONNECTED,
      PCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_17_UNCONNECTED,
      PCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_16_UNCONNECTED,
      PCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_15_UNCONNECTED,
      PCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_14_UNCONNECTED,
      PCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_13_UNCONNECTED,
      PCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_12_UNCONNECTED,
      PCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_11_UNCONNECTED,
      PCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_10_UNCONNECTED,
      PCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_9_UNCONNECTED,
      PCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_8_UNCONNECTED,
      PCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_7_UNCONNECTED,
      PCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_6_UNCONNECTED,
      PCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_5_UNCONNECTED,
      PCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_4_UNCONNECTED,
      PCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_3_UNCONNECTED,
      PCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_2_UNCONNECTED,
      PCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_1_UNCONNECTED,
      PCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_PCOUT_0_UNCONNECTED,
      ACOUT(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_29_UNCONNECTED,
      ACOUT(28) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_28_UNCONNECTED,
      ACOUT(27) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_27_UNCONNECTED,
      ACOUT(26) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_26_UNCONNECTED,
      ACOUT(25) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_25_UNCONNECTED,
      ACOUT(24) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_24_UNCONNECTED,
      ACOUT(23) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_23_UNCONNECTED,
      ACOUT(22) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_22_UNCONNECTED,
      ACOUT(21) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_21_UNCONNECTED,
      ACOUT(20) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_20_UNCONNECTED,
      ACOUT(19) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_19_UNCONNECTED,
      ACOUT(18) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_18_UNCONNECTED,
      ACOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_17_UNCONNECTED,
      ACOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_16_UNCONNECTED,
      ACOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_15_UNCONNECTED,
      ACOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_14_UNCONNECTED,
      ACOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_13_UNCONNECTED,
      ACOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_12_UNCONNECTED,
      ACOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_11_UNCONNECTED,
      ACOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_10_UNCONNECTED,
      ACOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_9_UNCONNECTED,
      ACOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_8_UNCONNECTED,
      ACOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_7_UNCONNECTED,
      ACOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_6_UNCONNECTED,
      ACOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_5_UNCONNECTED,
      ACOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_4_UNCONNECTED,
      ACOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_3_UNCONNECTED,
      ACOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_2_UNCONNECTED,
      ACOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_1_UNCONNECTED,
      ACOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_ACOUT_0_UNCONNECTED,
      OPMODE(6) => blk00000001_blk000001a2_sig00000592,
      OPMODE(5) => blk00000001_blk000001a2_sig00000592,
      OPMODE(4) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(3) => blk00000001_blk000001a2_sig00000592,
      OPMODE(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      OPMODE(1) => blk00000001_blk000001a2_sig00000592,
      OPMODE(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CARRYOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_3_UNCONNECTED,
      CARRYOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_2_UNCONNECTED,
      CARRYOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_1_UNCONNECTED,
      CARRYOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_CARRYOUT_0_UNCONNECTED,
      BCIN(17) => blk00000001_blk000001a2_sig00000592,
      BCIN(16) => blk00000001_blk000001a2_sig00000592,
      BCIN(15) => blk00000001_blk000001a2_sig00000592,
      BCIN(14) => blk00000001_blk000001a2_sig00000592,
      BCIN(13) => blk00000001_blk000001a2_sig00000592,
      BCIN(12) => blk00000001_blk000001a2_sig00000592,
      BCIN(11) => blk00000001_blk000001a2_sig00000592,
      BCIN(10) => blk00000001_blk000001a2_sig00000592,
      BCIN(9) => blk00000001_blk000001a2_sig00000592,
      BCIN(8) => blk00000001_blk000001a2_sig00000592,
      BCIN(7) => blk00000001_blk000001a2_sig00000592,
      BCIN(6) => blk00000001_blk000001a2_sig00000592,
      BCIN(5) => blk00000001_blk000001a2_sig00000592,
      BCIN(4) => blk00000001_blk000001a2_sig00000592,
      BCIN(3) => blk00000001_blk000001a2_sig00000592,
      BCIN(2) => blk00000001_blk000001a2_sig00000592,
      BCIN(1) => blk00000001_blk000001a2_sig00000592,
      BCIN(0) => blk00000001_blk000001a2_sig00000592,
      BCOUT(17) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_17_UNCONNECTED,
      BCOUT(16) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_16_UNCONNECTED,
      BCOUT(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_15_UNCONNECTED,
      BCOUT(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_14_UNCONNECTED,
      BCOUT(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_13_UNCONNECTED,
      BCOUT(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_12_UNCONNECTED,
      BCOUT(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_11_UNCONNECTED,
      BCOUT(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_10_UNCONNECTED,
      BCOUT(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_9_UNCONNECTED,
      BCOUT(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_8_UNCONNECTED,
      BCOUT(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_7_UNCONNECTED,
      BCOUT(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_6_UNCONNECTED,
      BCOUT(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_5_UNCONNECTED,
      BCOUT(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_4_UNCONNECTED,
      BCOUT(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_3_UNCONNECTED,
      BCOUT(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_2_UNCONNECTED,
      BCOUT(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_1_UNCONNECTED,
      BCOUT(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115d_BCOUT_0_UNCONNECTED,
      ACIN(29) => blk00000001_blk000001a2_sig00000592,
      ACIN(28) => blk00000001_blk000001a2_sig00000592,
      ACIN(27) => blk00000001_blk000001a2_sig00000592,
      ACIN(26) => blk00000001_blk000001a2_sig00000592,
      ACIN(25) => blk00000001_blk000001a2_sig00000592,
      ACIN(24) => blk00000001_blk000001a2_sig00000592,
      ACIN(23) => blk00000001_blk000001a2_sig00000592,
      ACIN(22) => blk00000001_blk000001a2_sig00000592,
      ACIN(21) => blk00000001_blk000001a2_sig00000592,
      ACIN(20) => blk00000001_blk000001a2_sig00000592,
      ACIN(19) => blk00000001_blk000001a2_sig00000592,
      ACIN(18) => blk00000001_blk000001a2_sig00000592,
      ACIN(17) => blk00000001_blk000001a2_sig00000592,
      ACIN(16) => blk00000001_blk000001a2_sig00000592,
      ACIN(15) => blk00000001_blk000001a2_sig00000592,
      ACIN(14) => blk00000001_blk000001a2_sig00000592,
      ACIN(13) => blk00000001_blk000001a2_sig00000592,
      ACIN(12) => blk00000001_blk000001a2_sig00000592,
      ACIN(11) => blk00000001_blk000001a2_sig00000592,
      ACIN(10) => blk00000001_blk000001a2_sig00000592,
      ACIN(9) => blk00000001_blk000001a2_sig00000592,
      ACIN(8) => blk00000001_blk000001a2_sig00000592,
      ACIN(7) => blk00000001_blk000001a2_sig00000592,
      ACIN(6) => blk00000001_blk000001a2_sig00000592,
      ACIN(5) => blk00000001_blk000001a2_sig00000592,
      ACIN(4) => blk00000001_blk000001a2_sig00000592,
      ACIN(3) => blk00000001_blk000001a2_sig00000592,
      ACIN(2) => blk00000001_blk000001a2_sig00000592,
      ACIN(1) => blk00000001_blk000001a2_sig00000592,
      ACIN(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001402,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001354
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115b : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001402,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk0000115b_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000115a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001401,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001353
    );
  blk00000001_blk000001a2_blk000001a3_blk00001159 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001401,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00001159_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00001158 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001400,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001351
    );
  blk00000001_blk000001a2_blk000001a3_blk00001157 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001400,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00001157_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00001156 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ff,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001232
    );
  blk00000001_blk000001a2_blk000001a3_blk00001155 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000124b,
      Q => blk00000001_blk000001a2_blk000001a3_sig000013ff,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00001155_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00001154 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013fe,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001352
    );
  blk00000001_blk000001a2_blk000001a3_blk00001153 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135d,
      Q => blk00000001_blk000001a2_blk000001a3_sig000013fe,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00001153_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00001152 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000009a,
      ENBWREN => blk00000001_sig0000009a,
      REGCEAREGCE => blk00000001_sig0000009a,
      REGCEB => blk00000001_sig0000009a,
      RSTRAMARSTRAM => blk00000001_blk000001a2_sig00000592,
      RSTRAMB => blk00000001_blk000001a2_sig00000592,
      RSTREGARSTREG => blk00000001_blk000001a2_sig00000592,
      RSTREGB => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(9) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011cd,
      ADDRARDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011cc,
      ADDRARDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011cb,
      ADDRARDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011ca,
      ADDRARDADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011c9,
      ADDRARDADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011cd,
      ADDRBWRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011cc,
      ADDRBWRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011cb,
      ADDRBWRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011ca,
      ADDRBWRADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011c9,
      ADDRBWRADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DIADI(15) => blk00000001_blk000001a2_sig00000592,
      DIADI(14) => blk00000001_blk000001a2_sig00000592,
      DIADI(13) => blk00000001_blk000001a2_sig00000592,
      DIADI(12) => blk00000001_blk000001a2_sig00000592,
      DIADI(11) => blk00000001_blk000001a2_sig00000592,
      DIADI(10) => blk00000001_blk000001a2_sig00000592,
      DIADI(9) => blk00000001_blk000001a2_sig00000592,
      DIADI(8) => blk00000001_blk000001a2_sig00000592,
      DIADI(7) => blk00000001_blk000001a2_sig00000592,
      DIADI(6) => blk00000001_blk000001a2_sig00000592,
      DIADI(5) => blk00000001_blk000001a2_sig00000592,
      DIADI(4) => blk00000001_blk000001a2_sig00000592,
      DIADI(3) => blk00000001_blk000001a2_sig00000592,
      DIADI(2) => blk00000001_blk000001a2_sig00000592,
      DIADI(1) => blk00000001_blk000001a2_sig00000592,
      DIADI(0) => blk00000001_blk000001a2_sig00000592,
      DIBDI(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => blk00000001_blk000001a2_sig00000592,
      DIPADIP(0) => blk00000001_blk000001a2_sig00000592,
      DIPBDIP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_blk000001a2_blk000001a3_sig000013d7,
      DOADO(14) => blk00000001_blk000001a2_blk000001a3_sig000013d6,
      DOADO(13) => blk00000001_blk000001a2_blk000001a3_sig000013d5,
      DOADO(12) => blk00000001_blk000001a2_blk000001a3_sig000013d4,
      DOADO(11) => blk00000001_blk000001a2_blk000001a3_sig000013d3,
      DOADO(10) => blk00000001_blk000001a2_blk000001a3_sig000013d2,
      DOADO(9) => blk00000001_blk000001a2_blk000001a3_sig000013d1,
      DOADO(8) => blk00000001_blk000001a2_blk000001a3_sig000013d0,
      DOADO(7) => blk00000001_blk000001a2_blk000001a3_sig000013cf,
      DOADO(6) => blk00000001_blk000001a2_blk000001a3_sig000013ce,
      DOADO(5) => blk00000001_blk000001a2_blk000001a3_sig000013cd,
      DOADO(4) => blk00000001_blk000001a2_blk000001a3_sig000013cc,
      DOADO(3) => blk00000001_blk000001a2_blk000001a3_sig000013cb,
      DOADO(2) => blk00000001_blk000001a2_blk000001a3_sig000013ca,
      DOADO(1) => blk00000001_blk000001a2_blk000001a3_sig000013c9,
      DOADO(0) => blk00000001_blk000001a2_blk000001a3_sig000013c8,
      DOBDO(15) => blk00000001_blk000001a2_blk000001a3_sig000013c6,
      DOBDO(14) => blk00000001_blk000001a2_blk000001a3_sig000013c5,
      DOBDO(13) => blk00000001_blk000001a2_blk000001a3_sig000013c4,
      DOBDO(12) => blk00000001_blk000001a2_blk000001a3_sig000013c3,
      DOBDO(11) => blk00000001_blk000001a2_blk000001a3_sig000013c2,
      DOBDO(10) => blk00000001_blk000001a2_blk000001a3_sig000013c1,
      DOBDO(9) => blk00000001_blk000001a2_blk000001a3_sig000013c0,
      DOBDO(8) => blk00000001_blk000001a2_blk000001a3_sig000013bf,
      DOBDO(7) => blk00000001_blk000001a2_blk000001a3_sig000013be,
      DOBDO(6) => blk00000001_blk000001a2_blk000001a3_sig000013bd,
      DOBDO(5) => blk00000001_blk000001a2_blk000001a3_sig000013bc,
      DOBDO(4) => blk00000001_blk000001a2_blk000001a3_sig000013bb,
      DOBDO(3) => blk00000001_blk000001a2_blk000001a3_sig000013ba,
      DOBDO(2) => blk00000001_blk000001a2_blk000001a3_sig000013b9,
      DOBDO(1) => blk00000001_blk000001a2_blk000001a3_sig000013b8,
      DOBDO(0) => blk00000001_blk000001a2_blk000001a3_sig000013b7,
      DOPADOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_blk000001a2_blk000001a3_sig000013d8,
      DOPBDOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001152_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_blk000001a2_blk000001a3_sig000013c7,
      WEA(1) => blk00000001_blk000001a2_sig00000592,
      WEA(0) => blk00000001_blk000001a2_sig00000592,
      WEBWE(3) => blk00000001_blk000001a2_sig00000592,
      WEBWE(2) => blk00000001_blk000001a2_sig00000592,
      WEBWE(1) => blk00000001_blk000001a2_sig00000592,
      WEBWE(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001151 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000009a,
      ENBWREN => blk00000001_sig0000009a,
      REGCEAREGCE => blk00000001_sig0000009a,
      REGCEB => blk00000001_sig0000009a,
      RSTRAMARSTRAM => blk00000001_blk000001a2_sig00000592,
      RSTRAMB => blk00000001_blk000001a2_sig00000592,
      RSTREGARSTREG => blk00000001_blk000001a2_sig00000592,
      RSTREGB => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(9) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011d2,
      ADDRARDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011d1,
      ADDRARDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011d0,
      ADDRARDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011cf,
      ADDRARDADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011ce,
      ADDRARDADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011d2,
      ADDRBWRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011d1,
      ADDRBWRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011d0,
      ADDRBWRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011cf,
      ADDRBWRADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011ce,
      ADDRBWRADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DIADI(15) => blk00000001_blk000001a2_sig00000592,
      DIADI(14) => blk00000001_blk000001a2_sig00000592,
      DIADI(13) => blk00000001_blk000001a2_sig00000592,
      DIADI(12) => blk00000001_blk000001a2_sig00000592,
      DIADI(11) => blk00000001_blk000001a2_sig00000592,
      DIADI(10) => blk00000001_blk000001a2_sig00000592,
      DIADI(9) => blk00000001_blk000001a2_sig00000592,
      DIADI(8) => blk00000001_blk000001a2_sig00000592,
      DIADI(7) => blk00000001_blk000001a2_sig00000592,
      DIADI(6) => blk00000001_blk000001a2_sig00000592,
      DIADI(5) => blk00000001_blk000001a2_sig00000592,
      DIADI(4) => blk00000001_blk000001a2_sig00000592,
      DIADI(3) => blk00000001_blk000001a2_sig00000592,
      DIADI(2) => blk00000001_blk000001a2_sig00000592,
      DIADI(1) => blk00000001_blk000001a2_sig00000592,
      DIADI(0) => blk00000001_blk000001a2_sig00000592,
      DIBDI(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => blk00000001_blk000001a2_sig00000592,
      DIPADIP(0) => blk00000001_blk000001a2_sig00000592,
      DIPBDIP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_blk000001a2_blk000001a3_sig000013b5,
      DOADO(14) => blk00000001_blk000001a2_blk000001a3_sig000013b4,
      DOADO(13) => blk00000001_blk000001a2_blk000001a3_sig000013b3,
      DOADO(12) => blk00000001_blk000001a2_blk000001a3_sig000013b2,
      DOADO(11) => blk00000001_blk000001a2_blk000001a3_sig000013b1,
      DOADO(10) => blk00000001_blk000001a2_blk000001a3_sig000013b0,
      DOADO(9) => blk00000001_blk000001a2_blk000001a3_sig000013af,
      DOADO(8) => blk00000001_blk000001a2_blk000001a3_sig000013ae,
      DOADO(7) => blk00000001_blk000001a2_blk000001a3_sig000013ad,
      DOADO(6) => blk00000001_blk000001a2_blk000001a3_sig000013ac,
      DOADO(5) => blk00000001_blk000001a2_blk000001a3_sig000013ab,
      DOADO(4) => blk00000001_blk000001a2_blk000001a3_sig000013aa,
      DOADO(3) => blk00000001_blk000001a2_blk000001a3_sig000013a9,
      DOADO(2) => blk00000001_blk000001a2_blk000001a3_sig000013a8,
      DOADO(1) => blk00000001_blk000001a2_blk000001a3_sig000013a7,
      DOADO(0) => blk00000001_blk000001a2_blk000001a3_sig000013a6,
      DOBDO(15) => blk00000001_blk000001a2_blk000001a3_sig000013a4,
      DOBDO(14) => blk00000001_blk000001a2_blk000001a3_sig000013a3,
      DOBDO(13) => blk00000001_blk000001a2_blk000001a3_sig000013a2,
      DOBDO(12) => blk00000001_blk000001a2_blk000001a3_sig000013a1,
      DOBDO(11) => blk00000001_blk000001a2_blk000001a3_sig000013a0,
      DOBDO(10) => blk00000001_blk000001a2_blk000001a3_sig0000139f,
      DOBDO(9) => blk00000001_blk000001a2_blk000001a3_sig0000139e,
      DOBDO(8) => blk00000001_blk000001a2_blk000001a3_sig0000139d,
      DOBDO(7) => blk00000001_blk000001a2_blk000001a3_sig0000139c,
      DOBDO(6) => blk00000001_blk000001a2_blk000001a3_sig0000139b,
      DOBDO(5) => blk00000001_blk000001a2_blk000001a3_sig0000139a,
      DOBDO(4) => blk00000001_blk000001a2_blk000001a3_sig00001399,
      DOBDO(3) => blk00000001_blk000001a2_blk000001a3_sig00001398,
      DOBDO(2) => blk00000001_blk000001a2_blk000001a3_sig00001397,
      DOBDO(1) => blk00000001_blk000001a2_blk000001a3_sig00001396,
      DOBDO(0) => blk00000001_blk000001a2_blk000001a3_sig00001395,
      DOPADOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_blk000001a2_blk000001a3_sig000013b6,
      DOPBDOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001151_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_blk000001a2_blk000001a3_sig000013a5,
      WEA(1) => blk00000001_blk000001a2_sig00000592,
      WEA(0) => blk00000001_blk000001a2_sig00000592,
      WEBWE(3) => blk00000001_blk000001a2_sig00000592,
      WEBWE(2) => blk00000001_blk000001a2_sig00000592,
      WEBWE(1) => blk00000001_blk000001a2_sig00000592,
      WEBWE(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk00001150 : RAMB18E1
    generic map(
      INITP_00 => X"0000000000000000000000000000000055555554000000000000000000000000",
      INIT_00 => X"7F627D8A7A7D764270E36A6E62F25A825134471D3C5730FC252818F90C8C0000",
      INIT_01 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_02 => X"0C8C18F9252830FC3C57471D51345A8262F26A6E70E376427A7D7D8A7F628000",
      INIT_03 => X"809E8276858389BE8F1D95929D0EA57EAECCB8E3C3A9CF04DAD8E707F3740000",
      INIT_A => X"00000",
      INIT_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      DOA_REG => 1,
      DOB_REG => 1,
      READ_WIDTH_A => 18,
      READ_WIDTH_B => 18,
      WRITE_WIDTH_A => 18,
      WRITE_WIDTH_B => 0,
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      RSTREG_PRIORITY_A => "RSTREG",
      RSTREG_PRIORITY_B => "RSTREG",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      SIM_COLLISION_CHECK => "ALL",
      INIT_FILE => "NONE"
    )
    port map (
      CLKARDCLK => aclk,
      CLKBWRCLK => aclk,
      ENARDEN => blk00000001_sig0000009a,
      ENBWREN => blk00000001_sig0000009a,
      REGCEAREGCE => blk00000001_sig0000009a,
      REGCEB => blk00000001_sig0000009a,
      RSTRAMARSTRAM => blk00000001_blk000001a2_sig00000592,
      RSTRAMB => blk00000001_blk000001a2_sig00000592,
      RSTREGARSTREG => blk00000001_blk000001a2_sig00000592,
      RSTREGB => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(9) => blk00000001_blk000001a2_sig00000592,
      ADDRARDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011d7,
      ADDRARDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011d6,
      ADDRARDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011d5,
      ADDRARDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011d4,
      ADDRARDADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011d3,
      ADDRARDADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRARDADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(13) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(12) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(11) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(10) => blk00000001_blk000001a2_sig00000592,
      ADDRBWRADDR(9) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000011d7,
      ADDRBWRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000011d6,
      ADDRBWRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000011d5,
      ADDRBWRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000011d4,
      ADDRBWRADDR(4) => blk00000001_blk000001a2_blk000001a3_sig000011d3,
      ADDRBWRADDR(3) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(2) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(1) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      ADDRBWRADDR(0) => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DIADI(15) => blk00000001_blk000001a2_sig00000592,
      DIADI(14) => blk00000001_blk000001a2_sig00000592,
      DIADI(13) => blk00000001_blk000001a2_sig00000592,
      DIADI(12) => blk00000001_blk000001a2_sig00000592,
      DIADI(11) => blk00000001_blk000001a2_sig00000592,
      DIADI(10) => blk00000001_blk000001a2_sig00000592,
      DIADI(9) => blk00000001_blk000001a2_sig00000592,
      DIADI(8) => blk00000001_blk000001a2_sig00000592,
      DIADI(7) => blk00000001_blk000001a2_sig00000592,
      DIADI(6) => blk00000001_blk000001a2_sig00000592,
      DIADI(5) => blk00000001_blk000001a2_sig00000592,
      DIADI(4) => blk00000001_blk000001a2_sig00000592,
      DIADI(3) => blk00000001_blk000001a2_sig00000592,
      DIADI(2) => blk00000001_blk000001a2_sig00000592,
      DIADI(1) => blk00000001_blk000001a2_sig00000592,
      DIADI(0) => blk00000001_blk000001a2_sig00000592,
      DIBDI(15) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_15_UNCONNECTED,
      DIBDI(14) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_14_UNCONNECTED,
      DIBDI(13) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_13_UNCONNECTED,
      DIBDI(12) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_12_UNCONNECTED,
      DIBDI(11) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_11_UNCONNECTED,
      DIBDI(10) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_10_UNCONNECTED,
      DIBDI(9) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_9_UNCONNECTED,
      DIBDI(8) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_8_UNCONNECTED,
      DIBDI(7) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_7_UNCONNECTED,
      DIBDI(6) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_6_UNCONNECTED,
      DIBDI(5) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_5_UNCONNECTED,
      DIBDI(4) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_4_UNCONNECTED,
      DIBDI(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_3_UNCONNECTED,
      DIBDI(2) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_2_UNCONNECTED,
      DIBDI(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_1_UNCONNECTED,
      DIBDI(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIBDI_0_UNCONNECTED,
      DIPADIP(1) => blk00000001_blk000001a2_sig00000592,
      DIPADIP(0) => blk00000001_blk000001a2_sig00000592,
      DIPBDIP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIPBDIP_1_UNCONNECTED,
      DIPBDIP(0) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DIPBDIP_0_UNCONNECTED,
      DOADO(15) => blk00000001_blk000001a2_blk000001a3_sig00001393,
      DOADO(14) => blk00000001_blk000001a2_blk000001a3_sig00001392,
      DOADO(13) => blk00000001_blk000001a2_blk000001a3_sig00001391,
      DOADO(12) => blk00000001_blk000001a2_blk000001a3_sig00001390,
      DOADO(11) => blk00000001_blk000001a2_blk000001a3_sig0000138f,
      DOADO(10) => blk00000001_blk000001a2_blk000001a3_sig0000138e,
      DOADO(9) => blk00000001_blk000001a2_blk000001a3_sig0000138d,
      DOADO(8) => blk00000001_blk000001a2_blk000001a3_sig0000138c,
      DOADO(7) => blk00000001_blk000001a2_blk000001a3_sig0000138b,
      DOADO(6) => blk00000001_blk000001a2_blk000001a3_sig0000138a,
      DOADO(5) => blk00000001_blk000001a2_blk000001a3_sig00001389,
      DOADO(4) => blk00000001_blk000001a2_blk000001a3_sig00001388,
      DOADO(3) => blk00000001_blk000001a2_blk000001a3_sig00001387,
      DOADO(2) => blk00000001_blk000001a2_blk000001a3_sig00001386,
      DOADO(1) => blk00000001_blk000001a2_blk000001a3_sig00001385,
      DOADO(0) => blk00000001_blk000001a2_blk000001a3_sig00001384,
      DOBDO(15) => blk00000001_blk000001a2_blk000001a3_sig00001382,
      DOBDO(14) => blk00000001_blk000001a2_blk000001a3_sig00001381,
      DOBDO(13) => blk00000001_blk000001a2_blk000001a3_sig00001380,
      DOBDO(12) => blk00000001_blk000001a2_blk000001a3_sig0000137f,
      DOBDO(11) => blk00000001_blk000001a2_blk000001a3_sig0000137e,
      DOBDO(10) => blk00000001_blk000001a2_blk000001a3_sig0000137d,
      DOBDO(9) => blk00000001_blk000001a2_blk000001a3_sig0000137c,
      DOBDO(8) => blk00000001_blk000001a2_blk000001a3_sig0000137b,
      DOBDO(7) => blk00000001_blk000001a2_blk000001a3_sig0000137a,
      DOBDO(6) => blk00000001_blk000001a2_blk000001a3_sig00001379,
      DOBDO(5) => blk00000001_blk000001a2_blk000001a3_sig00001378,
      DOBDO(4) => blk00000001_blk000001a2_blk000001a3_sig00001377,
      DOBDO(3) => blk00000001_blk000001a2_blk000001a3_sig00001376,
      DOBDO(2) => blk00000001_blk000001a2_blk000001a3_sig00001375,
      DOBDO(1) => blk00000001_blk000001a2_blk000001a3_sig00001374,
      DOBDO(0) => blk00000001_blk000001a2_blk000001a3_sig00001373,
      DOPADOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DOPADOP_1_UNCONNECTED,
      DOPADOP(0) => blk00000001_blk000001a2_blk000001a3_sig00001394,
      DOPBDOP(1) => NLW_blk00000001_blk000001a2_blk000001a3_blk00001150_DOPBDOP_1_UNCONNECTED,
      DOPBDOP(0) => blk00000001_blk000001a2_blk000001a3_sig00001383,
      WEA(1) => blk00000001_blk000001a2_sig00000592,
      WEA(0) => blk00000001_blk000001a2_sig00000592,
      WEBWE(3) => blk00000001_blk000001a2_sig00000592,
      WEBWE(2) => blk00000001_blk000001a2_sig00000592,
      WEBWE(1) => blk00000001_blk000001a2_sig00000592,
      WEBWE(0) => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114f : LUT5
    generic map(
      INIT => X"55551555"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012a2,
      I3 => blk00000001_sig0000009a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000012a1,
      O => blk00000001_blk000001a2_blk000001a3_sig000013fd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114e : LUT6
    generic map(
      INIT => X"4044444444444444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012a1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000012a5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000012a2,
      I5 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000013fc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114d : MUXF7
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000013fc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000013fd,
      S => blk00000001_blk000001a2_blk000001a3_sig0000126b,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114c : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig0000126a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001223
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114b : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001269,
      O => blk00000001_blk000001a2_blk000001a3_sig00001222
    );
  blk00000001_blk000001a2_blk000001a3_blk0000114a : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001268,
      O => blk00000001_blk000001a2_blk000001a3_sig00001221
    );
  blk00000001_blk000001a2_blk000001a3_blk00001149 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001267,
      O => blk00000001_blk000001a2_blk000001a3_sig00001220
    );
  blk00000001_blk000001a2_blk000001a3_blk00001148 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001266,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001147 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001265,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001146 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00000e27,
      O => blk00000001_blk000001a2_blk000001a3_sig00000df6
    );
  blk00000001_blk000001a2_blk000001a3_blk00001145 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00000d40,
      O => blk00000001_blk000001a2_blk000001a3_sig00000d83
    );
  blk00000001_blk000001a2_blk000001a3_blk00001144 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00000d40,
      O => blk00000001_blk000001a2_blk000001a3_sig00000d0f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001143 : LUT3
    generic map(
      INIT => X"FB"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000124b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011f6,
      I2 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig000011b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00001142 : LUT4
    generic map(
      INIT => X"1F0A"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001232,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124b,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00001141 : LUT4
    generic map(
      INIT => X"1F0A"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001249,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124a,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001140 : LUT6
    generic map(
      INIT => X"FFFFFFFF88880800"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_sig00000099,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      O => blk00000001_blk000001a2_blk000001a3_sig000012cd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113f : LUT5
    generic map(
      INIT => X"FFFF2000"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I2 => blk00000001_blk000001a2_sig00000753,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000012c3,
      O => blk00000001_blk000001a2_blk000001a3_sig000012be
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113e : LUT5
    generic map(
      INIT => X"FFFF8000"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I2 => blk00000001_blk000001a2_sig00000753,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001200,
      O => blk00000001_blk000001a2_blk000001a3_sig000012af
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113d : LUT5
    generic map(
      INIT => X"AAAA222A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012a6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001294
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113c : LUT4
    generic map(
      INIT => X"FF80"
    )
    port map (
      I0 => blk00000001_sig000000c7,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I3 => blk00000001_sig0000009b,
      O => blk00000001_blk000001a2_blk000001a3_sig00001278
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113b : LUT6
    generic map(
      INIT => X"AAAAFEAA00000000"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I4 => blk00000001_sig00000099,
      I5 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001299
    );
  blk00000001_blk000001a2_blk000001a3_blk0000113a : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001231,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00001139 : LUT6
    generic map(
      INIT => X"0454044404440444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00001138 : LUT5
    generic map(
      INIT => X"FFEAFF2A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000090d,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_sig00000097,
      I3 => blk00000001_sig00000099,
      I4 => blk00000001_sig00000098,
      O => blk00000001_blk000001a2_blk000001a3_sig000013ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00001137 : LUT6
    generic map(
      INIT => X"5410101010101010"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      I4 => blk00000001_blk000001a2_sig00000753,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00001136 : LUT6
    generic map(
      INIT => X"0111010100100000"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000124b,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000007fd,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090b,
      I5 => blk00000001_sig000000cb,
      O => blk00000001_blk000001a2_blk000001a3_sig000013ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00001135 : LUT5
    generic map(
      INIT => X"04540444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_sig00000753,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      O => blk00000001_blk000001a2_blk000001a3_sig000013ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00001134 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001257,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00001133 : LUT5
    generic map(
      INIT => X"51114000"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      I4 => blk00000001_sig000000c8,
      O => blk00000001_blk000001a2_blk000001a3_sig000013ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00001132 : LUT5
    generic map(
      INIT => X"04540444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a1,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000012a6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000129a,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00001131 : LUT6
    generic map(
      INIT => X"0454044404440444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000090b,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000007fb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007fa,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000990,
      O => blk00000001_blk000001a2_blk000001a3_sig000013ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00001130 : LUT5
    generic map(
      INIT => X"FFFF3A2A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000124e,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I4 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112f : LUT6
    generic map(
      INIT => X"0444044404540444"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig000000c7,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I4 => blk00000001_sig00000096,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000013fb,
      O => blk00000001_blk000001a2_blk000001a3_sig000013eb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112e : LUT4
    generic map(
      INIT => X"FF01"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001231,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      O => blk00000001_blk000001a2_blk000001a3_sig000013fb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112d : LUT6
    generic map(
      INIT => X"ECECEEECCCCCCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      I4 => blk00000001_sig00000099,
      I5 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012cc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112c : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012c2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012bd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112b : LUT5
    generic map(
      INIT => X"ECCCCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000124e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ae
    );
  blk00000001_blk000001a2_blk000001a3_blk0000112a : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001240,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001255,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001293
    );
  blk00000001_blk000001a2_blk000001a3_blk00001129 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig0000009c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001277
    );
  blk00000001_blk000001a2_blk000001a3_blk00001128 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012c1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00001127 : LUT5
    generic map(
      INIT => X"EAAAAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000124e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00001126 : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001254,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001292
    );
  blk00000001_blk000001a2_blk000001a3_blk00001125 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig0000009d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001276
    );
  blk00000001_blk000001a2_blk000001a3_blk00001124 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012c0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00001123 : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001253,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001291
    );
  blk00000001_blk000001a2_blk000001a3_blk00001122 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig0000009e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001275
    );
  blk00000001_blk000001a2_blk000001a3_blk00001121 : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001252,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001290
    );
  blk00000001_blk000001a2_blk000001a3_blk00001120 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig0000009f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001274
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111f : LUT6
    generic map(
      INIT => X"FFFFFFFFFFFFFFFE"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000013de,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000013e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000013fa,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000013f5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000013dd,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000013e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001098
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111e : LUT5
    generic map(
      INIT => X"FFFF7FFE"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009c0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c46,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c45,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000013df,
      O => blk00000001_blk000001a2_blk000001a3_sig000013fa
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111d : LUT6
    generic map(
      INIT => X"FF00FFCCFF0EFFCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I3 => blk00000001_sig00000099,
      I4 => blk00000001_sig0000009a,
      I5 => blk00000001_sig00000096,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111c : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001251,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111b : LUT6
    generic map(
      INIT => X"FFF4FFFEFFF5FFFF"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c56,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000013e3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000013e2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000013f9,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000013f8,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000111a : LUT4
    generic map(
      INIT => X"AAAB"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c50,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c4f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00001119 : LUT6
    generic map(
      INIT => X"1010101010101011"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c55,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c50,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00000c4f,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000c4e,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00001118 : LUT6
    generic map(
      INIT => X"FFF7FFF2FFFFFFFA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c4d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000013db,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000013dc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000013f6,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000013f7,
      O => blk00000001_blk000001a2_blk000001a3_sig000013dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00001117 : LUT6
    generic map(
      INIT => X"8000000088888888"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c4c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c51,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00000c52,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000c53,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001116 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c53,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c52,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c51,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00001115 : LUT5
    generic map(
      INIT => X"00E00000"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I3 => blk00000001_sig00000099,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig0000126b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001114 : LUT6
    generic map(
      INIT => X"ECECEEECCCCCCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      I4 => blk00000001_sig00000099,
      I5 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00001113 : LUT5
    generic map(
      INIT => X"ECCCCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000124e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00001112 : LUT5
    generic map(
      INIT => X"AEAAAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012bf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I3 => blk00000001_blk000001a2_sig00000753,
      I4 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00001111 : LUT4
    generic map(
      INIT => X"EAAA"
    )
    port map (
      I0 => blk00000001_sig000000a0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001256,
      I2 => blk00000001_sig000000c7,
      I3 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001273
    );
  blk00000001_blk000001a2_blk000001a3_blk00001110 : LUT6
    generic map(
      INIT => X"CCCCCCCCAAACCCCC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000123b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001250,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I5 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110f : LUT5
    generic map(
      INIT => X"FFFF7FFE"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009a0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c40,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000013e1,
      O => blk00000001_blk000001a2_blk000001a3_sig000013f5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110e : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013f4,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110d : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013f3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001231
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110c : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013f2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001230
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110b : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013f1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000122f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000110a : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013f0,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000122e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001109 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ef,
      Q => blk00000001_sig000000c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00001108 : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ee,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000090d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001107 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ed,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000090b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001106 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ec,
      Q => blk00000001_sig000000cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00001105 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013eb,
      Q => blk00000001_sig000000c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001104 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ea,
      Q => blk00000001_blk000001a2_sig00000753
    );
  blk00000001_blk000001a2_blk000001a3_blk00001103 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013e9,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00001102 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013e8,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000124b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001101 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000124a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001100 : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013e6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001247
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ff : FD
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000013e5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001248
    );
  blk00000001_blk000001a2_blk000001a3_blk000010fe : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c44,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c43,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e3
    );
  blk00000001_blk000001a2_blk000001a3_blk000010fd : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c4d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c4c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e2
    );
  blk00000001_blk000001a2_blk000001a3_blk000010fc : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c53,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c52,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e1
    );
  blk00000001_blk000001a2_blk000001a3_blk000010fb : LUT4
    generic map(
      INIT => X"5554"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c4a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c49,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013e0
    );
  blk00000001_blk000001a2_blk000001a3_blk000010fa : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c44,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c43,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013df
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f9 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c4a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c49,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013de
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f8 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c50,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c4f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      O => blk00000001_blk000001a2_blk000001a3_sig000013dc
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f7 : LUT4
    generic map(
      INIT => X"2AAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c56,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c55,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      O => blk00000001_blk000001a2_blk000001a3_sig000013db
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f6 : LUT4
    generic map(
      INIT => X"9996"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001200,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      O => blk00000001_blk000001a2_blk000001a3_sig00001318
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f5 : LUT4
    generic map(
      INIT => X"9996"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001302,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001304,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001301,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001303,
      O => blk00000001_blk000001a2_blk000001a3_sig00001317
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      O => blk00000001_blk000001a2_blk000001a3_sig00001316
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001301,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001303,
      O => blk00000001_blk000001a2_blk000001a3_sig00001315
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f2 : LUT3
    generic map(
      INIT => X"02"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000012f3
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f1 : LUT3
    generic map(
      INIT => X"01"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000012f2
    );
  blk00000001_blk000001a2_blk000001a3_blk000010f0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001306,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001305,
      O => blk00000001_blk000001a2_blk000001a3_sig000012f1
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ef : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130b,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ee
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ee : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ed
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ed : LUT4
    generic map(
      INIT => X"AA9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e9
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ec : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130b,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e7
    );
  blk00000001_blk000001a2_blk000001a3_blk000010eb : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130b,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e8
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ea : LUT4
    generic map(
      INIT => X"AA9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e6
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e9 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e4
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e8 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001309,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012e5
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e7 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001300,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012ff,
      O => blk00000001_blk000001a2_blk000001a3_sig000012eb
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001300,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ff,
      O => blk00000001_blk000001a2_blk000001a3_sig000012f0
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ff,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001300,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ea
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e4 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ff,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ec
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ff,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ef
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e2 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001258,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000125a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00001259,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ce
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e1 : LUT3
    generic map(
      INIT => X"40"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012a1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012a4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000124f
    );
  blk00000001_blk000001a2_blk000001a3_blk000010e0 : LUT6
    generic map(
      INIT => X"2000000000000000"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001251,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001250,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001252,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001253,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001254,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00001255,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128c
    );
  blk00000001_blk000001a2_blk000001a3_blk000010df : LUT6
    generic map(
      INIT => X"2000000000000000"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001250,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001251,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001252,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001253,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001254,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00001255,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128d
    );
  blk00000001_blk000001a2_blk000001a3_blk000010de : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig00000097,
      O => blk00000001_blk000001a2_blk000001a3_sig0000122a
    );
  blk00000001_blk000001a2_blk000001a3_blk000010dd : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig000000c7,
      I1 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001229
    );
  blk00000001_blk000001a2_blk000001a3_blk000010dc : LUT3
    generic map(
      INIT => X"80"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I2 => blk00000001_blk000001a2_sig00000753,
      O => blk00000001_blk000001a2_blk000001a3_sig000011f9
    );
  blk00000001_blk000001a2_blk000001a3_blk000010db : LUT3
    generic map(
      INIT => X"40"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001247,
      I1 => blk00000001_sig0000009a,
      I2 => blk00000001_blk000001a2_sig00000753,
      O => blk00000001_blk000001a2_blk000001a3_sig00001227
    );
  blk00000001_blk000001a2_blk000001a3_blk000010da : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_sig000000c7,
      O => blk00000001_blk000001a2_blk000001a3_sig00001226
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d9 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000124b,
      O => blk00000001_blk000001a2_blk000001a3_sig000007f9
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d8 : LUT2
    generic map(
      INIT => X"E"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000124a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001225
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d7 : LUT4
    generic map(
      INIT => X"EEEF"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I1 => blk00000001_sig000000c7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001239,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000124c,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121d
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001209,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001203
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d5 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001204
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d4 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001205
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d3 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001206
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d2 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001207
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      O => blk00000001_blk000001a2_blk000001a3_sig00001208
    );
  blk00000001_blk000001a2_blk000001a3_blk000010d0 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001237,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001238,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121a
    );
  blk00000001_blk000001a2_blk000001a3_blk000010cf : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001238,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001237,
      O => blk00000001_blk000001a2_blk000001a3_sig00001219
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ce : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001238,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001237,
      O => blk00000001_blk000001a2_blk000001a3_sig00001218
    );
  blk00000001_blk000001a2_blk000001a3_blk000010cd : LUT2
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001238,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001237,
      O => blk00000001_blk000001a2_blk000001a3_sig00001217
    );
  blk00000001_blk000001a2_blk000001a3_blk000010cc : LUT6
    generic map(
      INIT => X"1010101010101000"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I1 => blk00000001_sig00000099,
      I2 => blk00000001_sig00000096,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00001231,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      O => blk00000001_blk000001a2_blk000001a3_sig000011fc
    );
  blk00000001_blk000001a2_blk000001a3_blk000010cb : LUT4
    generic map(
      INIT => X"00E0"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001230,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001248,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000122e,
      I3 => blk00000001_sig00000099,
      O => blk00000001_blk000001a2_blk000001a3_sig00001224
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ca : LUT5
    generic map(
      INIT => X"FF808080"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      I2 => blk00000001_blk000001a2_sig00000753,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000124f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121b
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c9 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      O => blk00000001_blk000001a2_blk000001a3_sig0000121c
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c8 : LUT4
    generic map(
      INIT => X"AA20"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig00000099,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000007fc,
      O => blk00000001_blk000001a2_blk000001a3_sig00001228
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c7 : LUT2
    generic map(
      INIT => X"4"
    )
    port map (
      I0 => blk00000001_sig00000099,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      O => blk00000001_blk000001a2_blk000001a3_sig000011fb
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c6 : LUT6
    generic map(
      INIT => X"56A9A9566A95956A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001212,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001211,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000122c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig00001210,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000122b,
      O => blk00000001_blk000001a2_blk000001a3_sig00001215
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c5 : LUT6
    generic map(
      INIT => X"56A9A9566A95956A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000120d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000120c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000120e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00001209,
      O => blk00000001_blk000001a2_blk000001a3_sig00001213
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c4 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000122b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001211,
      O => blk00000001_blk000001a2_blk000001a3_sig00001216
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c3 : LUT3
    generic map(
      INIT => X"96"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001209,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000120d,
      O => blk00000001_blk000001a2_blk000001a3_sig00001214
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c2 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011ea,
      O => blk00000001_blk000001a2_blk000001a3_sig000007ff
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011ed,
      I1 => blk00000001_sig0000009a,
      O => blk00000001_blk000001a2_blk000001a3_sig000007f6
    );
  blk00000001_blk000001a2_blk000001a3_blk000010c0 : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001236,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000011b2
    );
  blk00000001_blk000001a2_blk000001a3_blk000010bf : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001235,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000011b1
    );
  blk00000001_blk000001a2_blk000001a3_blk000010be : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001234,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000011b0
    );
  blk00000001_blk000001a2_blk000001a3_blk000010bd : LUT4
    generic map(
      INIT => X"D580"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001233,
      I2 => blk00000001_sig0000009a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ee,
      O => blk00000001_blk000001a2_blk000001a3_sig000011af
    );
  blk00000001_blk000001a2_blk000001a3_blk000010bc : LUT3
    generic map(
      INIT => X"4E"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      O => blk00000001_blk000001a2_blk000001a3_sig000010df
    );
  blk00000001_blk000001a2_blk000001a3_blk000010bb : LUT3
    generic map(
      INIT => X"1B"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      O => blk00000001_blk000001a2_blk000001a3_sig000010de
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ba : LUT3
    generic map(
      INIT => X"A9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      O => blk00000001_blk000001a2_blk000001a3_sig000010dd
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b9 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      O => blk00000001_blk000001a2_blk000001a3_sig000010dc
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b8 : LUT4
    generic map(
      INIT => X"78D8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000809,
      O => blk00000001_blk000001a2_blk000001a3_sig000010e0
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b7 : LUT4
    generic map(
      INIT => X"8D87"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000809,
      O => blk00000001_blk000001a2_blk000001a3_sig000010db
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b6 : LUT4
    generic map(
      INIT => X"D272"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000809,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d9
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b5 : LUT4
    generic map(
      INIT => X"272D"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000007f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000007e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007ea,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000809,
      O => blk00000001_blk000001a2_blk000001a3_sig000010da
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b4 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b20,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b34,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108d
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b3 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b33,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108c
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b2 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b32,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108b
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b1 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b31,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108a
    );
  blk00000001_blk000001a2_blk000001a3_blk000010b0 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b30,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001089
    );
  blk00000001_blk000001a2_blk000001a3_blk000010af : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001088
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ae : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001087
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ad : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b19,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001086
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ac : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001097
    );
  blk00000001_blk000001a2_blk000001a3_blk000010ab : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b29,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001096
    );
  blk00000001_blk000001a2_blk000001a3_blk000010aa : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b28,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001095
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a9 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b27,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001094
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a8 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b26,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001093
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a7 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b25,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001092
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a6 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b24,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001091
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a5 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b23,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001090
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a4 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b22,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b36,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108f
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a3 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b21,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b35,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000108e
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a2 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b18,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001085
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a1 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b17,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001084
    );
  blk00000001_blk000001a2_blk000001a3_blk000010a0 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b34,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001079
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109f : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b33,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001078
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109e : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b32,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001077
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109d : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b31,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001076
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109c : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b30,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001075
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109b : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001074
    );
  blk00000001_blk000001a2_blk000001a3_blk0000109a : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001073
    );
  blk00000001_blk000001a2_blk000001a3_blk00001099 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001072
    );
  blk00000001_blk000001a2_blk000001a3_blk00001098 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001083
    );
  blk00000001_blk000001a2_blk000001a3_blk00001097 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001082
    );
  blk00000001_blk000001a2_blk000001a3_blk00001096 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001081
    );
  blk00000001_blk000001a2_blk000001a3_blk00001095 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001080
    );
  blk00000001_blk000001a2_blk000001a3_blk00001094 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001093 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b39,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001092 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b38,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001091 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b37,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001090 : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b36,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108f : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b35,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000107a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108e : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001071
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108d : LUT3
    generic map(
      INIT => X"AC"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_sig00001070
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108c : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_sig00000097,
      O => blk00000001_blk000001a2_blk000001a3_sig0000090c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000809,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000090a,
      O => blk00000001_blk000001a2_blk000001a3_sig00000802
    );
  blk00000001_blk000001a2_blk000001a3_blk0000108a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013da,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00001089 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00001088 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001201,
      Q => blk00000001_blk000001a2_blk000001a3_sig000013da
    );
  blk00000001_blk000001a2_blk000001a3_blk00001087 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001202,
      Q => blk00000001_blk000001a2_blk000001a3_sig000013d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00001086 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e49
    );
  blk00000001_blk000001a2_blk000001a3_blk00001085 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001084 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ca,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001083 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013cb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001082 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013cc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001081 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013cd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001080 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ce,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e4f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013cf,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e50
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e51
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e52
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e53
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e54
    );
  blk00000001_blk000001a2_blk000001a3_blk0000107a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e55
    );
  blk00000001_blk000001a2_blk000001a3_blk00001079 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e56
    );
  blk00000001_blk000001a2_blk000001a3_blk00001078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e57
    );
  blk00000001_blk000001a2_blk000001a3_blk00001077 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e58
    );
  blk00000001_blk000001a2_blk000001a3_blk00001076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013d8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e59
    );
  blk00000001_blk000001a2_blk000001a3_blk00001075 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001074 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001073 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ba,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001071 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013bb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013bc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e5f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013bd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e60
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013be,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e61
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013bf,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e62
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e63
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e64
    );
  blk00000001_blk000001a2_blk000001a3_blk0000106a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e65
    );
  blk00000001_blk000001a2_blk000001a3_blk00001069 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e66
    );
  blk00000001_blk000001a2_blk000001a3_blk00001068 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e67
    );
  blk00000001_blk000001a2_blk000001a3_blk00001067 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e68
    );
  blk00000001_blk000001a2_blk000001a3_blk00001066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e69
    );
  blk00000001_blk000001a2_blk000001a3_blk00001065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013c7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e6a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd4
    );
  blk00000001_blk000001a2_blk000001a3_blk00001063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd5
    );
  blk00000001_blk000001a2_blk000001a3_blk00001062 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd6
    );
  blk00000001_blk000001a2_blk000001a3_blk00001061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013aa,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ab,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ac,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dda
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ad,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ddb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013ae,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ddc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013af,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ddd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000105a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dde
    );
  blk00000001_blk000001a2_blk000001a3_blk00001059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ddf
    );
  blk00000001_blk000001a2_blk000001a3_blk00001058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de0
    );
  blk00000001_blk000001a2_blk000001a3_blk00001057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de1
    );
  blk00000001_blk000001a2_blk000001a3_blk00001056 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de2
    );
  blk00000001_blk000001a2_blk000001a3_blk00001055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de3
    );
  blk00000001_blk000001a2_blk000001a3_blk00001054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013b6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de4
    );
  blk00000001_blk000001a2_blk000001a3_blk00001053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001395,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de5
    );
  blk00000001_blk000001a2_blk000001a3_blk00001052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001396,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de6
    );
  blk00000001_blk000001a2_blk000001a3_blk00001051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001397,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001050 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001398,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001399,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000de9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dea
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000deb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dec
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ded
    );
  blk00000001_blk000001a2_blk000001a3_blk0000104a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dee
    );
  blk00000001_blk000001a2_blk000001a3_blk00001049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000139f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000def
    );
  blk00000001_blk000001a2_blk000001a3_blk00001048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df0
    );
  blk00000001_blk000001a2_blk000001a3_blk00001047 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df1
    );
  blk00000001_blk000001a2_blk000001a3_blk00001046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df2
    );
  blk00000001_blk000001a2_blk000001a3_blk00001045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df3
    );
  blk00000001_blk000001a2_blk000001a3_blk00001044 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df4
    );
  blk00000001_blk000001a2_blk000001a3_blk00001043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000013a5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000df5
    );
  blk00000001_blk000001a2_blk000001a3_blk00001042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001384,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d61
    );
  blk00000001_blk000001a2_blk000001a3_blk00001041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001385,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d62
    );
  blk00000001_blk000001a2_blk000001a3_blk00001040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001386,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d63
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001387,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d64
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001388,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d65
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001389,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d66
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d67
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d68
    );
  blk00000001_blk000001a2_blk000001a3_blk0000103a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d69
    );
  blk00000001_blk000001a2_blk000001a3_blk00001039 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001038 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001037 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000138f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001036 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001390,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001035 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001391,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001034 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001392,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d6f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001033 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001393,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d70
    );
  blk00000001_blk000001a2_blk000001a3_blk00001032 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001394,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d71
    );
  blk00000001_blk000001a2_blk000001a3_blk00001031 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001373,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d72
    );
  blk00000001_blk000001a2_blk000001a3_blk00001030 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001374,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d73
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001375,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d74
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001376,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d75
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001377,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d76
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001378,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d77
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001379,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d78
    );
  blk00000001_blk000001a2_blk000001a3_blk0000102a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d79
    );
  blk00000001_blk000001a2_blk000001a3_blk00001029 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7a
    );
  blk00000001_blk000001a2_blk000001a3_blk00001028 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001027 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001026 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001025 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000137f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001024 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001380,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d7f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001023 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001381,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d80
    );
  blk00000001_blk000001a2_blk000001a3_blk00001022 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001382,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d81
    );
  blk00000001_blk000001a2_blk000001a3_blk00001021 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001383,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d82
    );
  blk00000001_blk000001a2_blk000001a3_blk00001020 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001372,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001371,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001370,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011de,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001372
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011df,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001371
    );
  blk00000001_blk000001a2_blk000001a3_blk0000101a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001370
    );
  blk00000001_blk000001a2_blk000001a3_blk00001019 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136f
    );
  blk00000001_blk000001a2_blk000001a3_blk00001018 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00001017 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011be
    );
  blk00000001_blk000001a2_blk000001a3_blk00001016 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00001015 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00001014 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136e
    );
  blk00000001_blk000001a2_blk000001a3_blk00001013 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e2,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136d
    );
  blk00000001_blk000001a2_blk000001a3_blk00001012 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e3,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136c
    );
  blk00000001_blk000001a2_blk000001a3_blk00001011 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e4,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136b
    );
  blk00000001_blk000001a2_blk000001a3_blk00001010 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000136a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001369,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ba
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001368,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011bb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001367,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011bc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011de,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000136a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001369
    );
  blk00000001_blk000001a2_blk000001a3_blk0000100a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001368
    );
  blk00000001_blk000001a2_blk000001a3_blk00001009 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001367
    );
  blk00000001_blk000001a2_blk000001a3_blk00001008 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001366,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00001007 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001365,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00001006 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001364,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00001005 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001363,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00001004 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001366
    );
  blk00000001_blk000001a2_blk000001a3_blk00001003 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001365
    );
  blk00000001_blk000001a2_blk000001a3_blk00001002 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001364
    );
  blk00000001_blk000001a2_blk000001a3_blk00001001 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011e9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001363
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001362,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000135e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001361,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000135d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001360,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000135c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000feb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000135b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fea : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011f2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011f4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ef,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000011f0,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001362
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe9 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011f1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011f3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ef,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000011f0,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001361
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe8 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011f2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ef,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000011f0,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001360
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe7 : LUT6
    generic map(
      INIT => X"00000000F0F0CCAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011f1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000011ef,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000011f0,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000135f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001354,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001353,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001352,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001351,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fe0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001354,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fdf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001353,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fde : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001352,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fdd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001351,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fdc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000135a,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fdb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001359,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011cd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fda : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001358,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011cc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001357,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001356,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001355,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001350,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001349
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134f,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000134a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134e,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000134b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134d,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000134c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001209,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001209,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001350
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120a,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000134f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fd0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120b,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000134e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fcf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120c,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000134d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fce : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120d,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fce_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fcd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000120e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000120e,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fcd_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fcc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001349,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134a,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134b,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011da
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000134c,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011db
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001348,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011dc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001347,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001306,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001300,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001348
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f0,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001347
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001346,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001345,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007db
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011de,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fc2_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011df,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001346
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fc0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fc0_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fbf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001345
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fbe : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001344,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fbd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001343,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007cd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fbc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001342,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007cc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fbb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001341,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fba : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011c1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001344
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011c2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001343
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011c3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001342
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011c4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001341
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001340,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007df
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fb4_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001340
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000fb2_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fb0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000faf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fac : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011bd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fab : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011be,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000faa : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011bf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011c0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000133a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007de
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001339,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001338,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007dc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001337,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011de,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig0000133a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001339
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001338
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001337
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fa0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001336,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001335,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001334,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001333,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011b9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001336
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011ba,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001335
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f9a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011bb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001334
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f99 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011bc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001333
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f98 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001332,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f97 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001331,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f96 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001330,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f95 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f94 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001332
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f93 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001331
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f92 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig00001330
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f91 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011e9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011ec,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f90 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007da
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011b5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011b6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f8a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011b7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f89 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011b8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000011c8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f88 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000132a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f87 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001329,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f86 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012fa,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f86_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f85 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ef,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000132a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f84 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f8,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f84_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f83 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f4,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001329
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f82 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001328,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f81 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001327,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f80 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012fa,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f80_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012ee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012eb,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001328
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f8,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f7e_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012ed,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001327
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001326,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001325,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f7a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001324,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f79 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001323,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f78 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012fa,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001326
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f77 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ec,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001325
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f76 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f8,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001324
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f75 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e4,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001323
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f74 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001322,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011de
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f73 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001321,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011df
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f72 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001320,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f71 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f70 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012fa,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001322
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012ea,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001321
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000012f8,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001320
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012e6,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000131f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f6a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012fc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f69 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012fb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f68 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001311,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001307,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001311,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000130c,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000130d,
      O => blk00000001_blk000001a2_blk000001a3_sig0000131e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f67 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001310,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001308,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001310,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000130c,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000130d,
      O => blk00000001_blk000001a2_blk000001a3_sig0000131d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f66 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001307,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000130f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130f,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000130c,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000130d,
      O => blk00000001_blk000001a2_blk000001a3_sig0000131c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f65 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001308,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000130e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000130e,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000130c,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000130d,
      O => blk00000001_blk000001a2_blk000001a3_sig0000131b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f50 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000131a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001306
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001319,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001305
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001308,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000131a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001307,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001319
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001318,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001307
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001317,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012ff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f4a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001316,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001308
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f49 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001315,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001300
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f48 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001314,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001309
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f47 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011f8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001314
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f46 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001313,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f45 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001312,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f44 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000012f2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001313
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f43 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000012f3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001312
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fe,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001310
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001200,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001311
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000130d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001301,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001302,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001303,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012fb,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f38 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012fc,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f37 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012fd,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f36 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012fe,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f35 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012e3,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f34 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012e2,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f33 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012e1,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f32 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012e0,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f31 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012df,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f30 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012de,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2f : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001203,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001204,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001205,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2c : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001206,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012e0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2b : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001207,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012df
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f2a : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001208,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012de
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f29 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012dd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f28 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012dc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f27 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f26 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012dc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012db,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012da,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f10_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0f : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012db
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0e : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012da
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0d : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f0a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f09 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f08 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f07 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fe,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f06 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f05 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001200,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f04 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f03 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f02 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f01 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f00 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000120f,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eff : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001210,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000efe : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001211,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000efd : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001212,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000efc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012d0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000efb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012cf,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000efa : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011dc,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ef9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_sig00000592,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011dd,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001228,
      D => blk00000001_blk000001a2_blk000001a3_sig000012ce,
      R => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001228,
      D => blk00000001_blk000001a2_blk000001a3_sig000012ca,
      R => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001228,
      D => blk00000001_blk000001a2_blk000001a3_sig000012c9,
      R => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001228,
      D => blk00000001_blk000001a2_blk000001a3_sig000012c8,
      R => blk00000001_blk000001a2_blk000001a3_sig0000122f,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb0 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012c2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012c3,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_sig00000592,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eaf : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012bf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012c0,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000012c1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eae : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig000012c4,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig000012c7,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ead : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig000012c6,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eac : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig000012c5,
      LI => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b9,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000124d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eaa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig0000124d,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007fc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ea9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b8,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012c3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ea8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b7,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012c2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ea7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b6,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012c1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ea6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b5,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ea5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001227,
      D => blk00000001_blk000001a2_blk000001a3_sig000012b4,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e97 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001200,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_sig00000592,
      I5 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e96 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000011fd,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000011fe,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000011ff,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e95 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig000012b0,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig000012b3,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e94 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig000012b2,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e93 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig000012b1,
      LI => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e92 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      D => blk00000001_blk000001a2_blk000001a3_sig000012ab,
      R => blk00000001_blk000001a2_blk000001a3_sig00001226,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000124e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e91 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      D => blk00000001_blk000001a2_blk000001a3_sig000012aa,
      R => blk00000001_blk000001a2_blk000001a3_sig00001226,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001200
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e90 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a9,
      R => blk00000001_blk000001a2_blk000001a3_sig00001226,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e8f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a8,
      R => blk00000001_blk000001a2_blk000001a3_sig00001226,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e8e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a7,
      R => blk00000001_blk000001a2_blk000001a3_sig00001226,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e77 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001224,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e76 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a3,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e75 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000129b,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig000000ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e74 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000129c,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e73 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000129d,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e72 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000129e,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e71 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000129f,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e70 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a0,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000129f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000012a1,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6e : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001287,
      S => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001286,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001255
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001285,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001254
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001284,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001253
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e6a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001283,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001252
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e69 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001282,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001251
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e68 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001299,
      D => blk00000001_blk000001a2_blk000001a3_sig00001281,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001250
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e67 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000127e,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e66 : FD
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000127d,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e65 : LUT3
    generic map(
      INIT => X"8A"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012a5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001298
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e64 : LUT3
    generic map(
      INIT => X"8A"
    )
    port map (
      I0 => blk00000001_sig0000009a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000012a5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001297
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e63 : LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001224,
      I3 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001296
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e62 : LUT4
    generic map(
      INIT => X"0001"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001224,
      I3 => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001295
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e61 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000127f,
      DI => blk00000001_blk000001a2_blk000001a3_sig000012a5,
      S => blk00000001_blk000001a2_blk000001a3_sig00001298,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e60 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00001280,
      DI => blk00000001_blk000001a2_blk000001a3_sig000012a4,
      S => blk00000001_blk000001a2_blk000001a3_sig00001297,
      O => blk00000001_blk000001a2_blk000001a3_sig0000128a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000128b,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig00001296,
      O => blk00000001_blk000001a2_blk000001a3_sig00001289
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000128a,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig00001295,
      O => blk00000001_blk000001a2_blk000001a3_sig00001288
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig0000128d,
      O => blk00000001_blk000001a2_blk000001a3_sig00001280
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig0000128c,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00001289,
      LI => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e5a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00001288,
      LI => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e46 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig0000009d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_sig0000009c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I4 => blk00000001_sig0000009b,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e45 : LUT6
    generic map(
      INIT => X"9009000000009009"
    )
    port map (
      I0 => blk00000001_sig000000a0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      I2 => blk00000001_sig0000009f,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_sig0000009e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e44 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00001279,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig0000127c,
      O => blk00000001_blk000001a2_blk000001a3_sig0000127a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e43 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig00000801,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_sig0000127b,
      O => blk00000001_blk000001a2_blk000001a3_sig00001279
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e42 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000127a,
      LI => blk00000001_blk000001a2_sig00000592,
      O => blk00000001_blk000001a2_blk000001a3_sig00001272
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e41 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig00001272,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001257
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e40 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig00001257,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001256
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig00001271,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig0000009b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig00001270,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig0000009c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig0000126f,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig0000009d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig0000126e,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig0000009e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig0000126d,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig0000009f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e3a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig00001229,
      D => blk00000001_blk000001a2_blk000001a3_sig0000126c,
      R => blk00000001_sig00000099,
      Q => blk00000001_sig000000a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e39 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig00000063,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001265
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e38 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig00000062,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001266
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e37 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig00000061,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001267
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e36 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig00000060,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001268
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e35 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig0000005f,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001269
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e34 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000122a,
      D => blk00000001_sig0000005e,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000126a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e33 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001241
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e32 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001242
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e31 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00001220,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001243
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e30 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00001221,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001244
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00001222,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001245
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00001223,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001246
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000800
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121b,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001217,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001233
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e2a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001218,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001234
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e29 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001235
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e28 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001219,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001236
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e27 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001225,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e26 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000121c,
      S => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000122d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e25 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001241,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e24 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001242,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e23 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001243,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e22 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001244,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e21 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001245,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000123f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e20 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001246,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001240
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig0000009c,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig0000009b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001210
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig0000009e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001211
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig0000009d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001212
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000012a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e1a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig000000a0,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000122b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e19 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_sig0000009f,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000122c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e18 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000124c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001239
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e17 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001250,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001209
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e16 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001251,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e15 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001252,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e14 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001253,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e13 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001254,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e12 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001255,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000120e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e11 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001216,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001237
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e10 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001215,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001238
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001214,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001201
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001213,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001202
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001264
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001263
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001262
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e0a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001261
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e09 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001260
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e08 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e07 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e06 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e05 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e04 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e03 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000125a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e02 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001259
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e01 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000801,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001258
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e00 : FDSE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011b3,
      S => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011af,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dfe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011b0,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dfd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011b1,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dfc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011b2,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dfb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fc,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d50 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ae,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ad,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008fb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ac,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008fc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011ab,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011aa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d4a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000900
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d49 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000901
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d48 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000902
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d47 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000903
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d46 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000904
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d45 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000905
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d44 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000906
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d43 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000907
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d42 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011a0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000908
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d41 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000909
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d40 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000950,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000951,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000952,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000953,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000954,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000955,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d3a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000956,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d39 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000957,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d38 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000958,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d37 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000959,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d36 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d35 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d34 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a53,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d33 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d32 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a55,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig000011a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d31 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000095f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a56,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d30 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000119a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001199,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d2a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001198,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d29 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001197,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d28 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001196,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d27 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001195,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d26 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001194,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d25 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001193,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d24 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001192,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d23 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001191,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d22 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001190,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d21 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d20 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000910,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000911,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000912,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000913,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000914,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000119a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000915,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001199
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d1a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000916,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001198
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d19 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000917,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001197
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d18 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000918,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001196
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d17 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000919,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001195
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d16 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001194
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d15 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001193
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d14 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001192
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d13 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001191
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d12 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001190
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d11 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000091f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008da
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008db
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008dc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000118a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008de
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001189,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008df
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d0a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001188,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d09 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001187,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d08 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001186,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d07 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001185,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d06 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001184,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d05 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001183,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d04 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001182,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d03 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001181,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d02 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001180,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d01 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008e9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d00 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000960,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cff : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000961,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cfe : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000962,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cfd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000963,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cfc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000964,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000118a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cfb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000965,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001189
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cfa : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000966,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001188
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000967,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001187
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000968,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001186
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000969,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001185
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001184
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001183
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a53,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001182
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001181
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a55,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001180
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000096f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a56,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cf0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008cc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ced : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008cd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000117a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ceb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001179,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001178,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001177,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001176,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001175,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001174,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001173,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001172,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001171,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001170,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ce0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000920,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cdf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000921,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cde : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000922,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cdd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000923,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cdc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000924,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000117a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cdb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000925,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001179
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cda : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000926,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001178
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000927,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001177
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000928,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001176
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000929,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001175
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001174
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001173
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001172
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001171
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001170
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000092f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cd0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ccf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ccd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ccc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000116a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008be
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ccb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001169,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001168,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001167,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001166,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001165,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001164,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001163,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001162,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001161,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001160,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cc0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000970,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cbf : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000971,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cbe : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000972,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cbd : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000973,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cbc : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000974,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000116a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cbb : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000975,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001169
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cba : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000976,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001168
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb9 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000977,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001167
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb8 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000978,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001166
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb7 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000979,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001165
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb6 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001164
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb5 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001163
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb4 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a53,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001162
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb3 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001161
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb2 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a55,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001160
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb1 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000097f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a56,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cb0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000caf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000115a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000cab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001159,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000caa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001158,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001157,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001156,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001155,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001154,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001153,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001152,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001151,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001150,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ca0 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000930,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000931,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000932,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000933,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000934,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000115a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000935,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001159
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c9a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000936,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001158
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c99 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000937,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001157
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c98 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000938,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001156
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c97 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000939,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001155
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c96 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001154
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c95 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001153
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c94 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001152
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c93 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001151
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c92 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001150
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c91 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000093f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c90 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000114a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001149,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000089f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c8a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001148,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c89 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001147,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c88 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001146,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c87 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001145,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c86 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001144,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c85 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001143,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c84 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001142,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c83 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001141,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c82 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001140,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c81 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000008a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c80 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000980,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000981,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000982,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000983,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000984,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000114a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000985,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001149
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c7a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000986,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001148
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c79 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000987,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001147
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c78 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000988,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001146
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c77 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000989,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001145
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c76 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001144
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c75 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001143
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c74 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a53,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001142
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c73 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a54,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001141
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c72 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a55,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001140
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c71 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000098f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a56,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c70 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000113a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001139,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000088f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c6a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001138,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000890
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c69 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001137,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000891
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c68 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001136,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000892
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c67 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001135,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000893
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c66 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001134,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000894
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c65 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001133,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000895
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c64 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001132,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000896
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c63 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001131,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000897
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c62 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001130,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000898
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c61 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000112f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000899
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c60 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000940,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5f : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000941,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5e : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000942,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5d : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000943,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5c : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000944,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000113a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5b : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000945,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001139
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c5a : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000946,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001138
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c59 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000947,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001137
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c58 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000948,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001136
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c57 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000949,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001135
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c56 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001134
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c55 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001133
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c54 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001132
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c53 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001131
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c52 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig00001130
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c51 : LUT3
    generic map(
      INIT => X"CA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000094f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000a46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000007f5,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c4a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000112a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000090f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c49 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001129,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000090e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c48 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000804,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000806,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000808,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c47 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000803,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000805,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000807,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c46 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c45 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_sig00000592,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ef,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007ee,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c44 : MUXF7
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000112e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000112c,
      S => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      O => blk00000001_blk000001a2_blk000001a3_sig0000112a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c43 : MUXF7
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000112d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000112b,
      S => blk00000001_blk000001a2_blk000001a3_sig000007ed,
      O => blk00000001_blk000001a2_blk000001a3_sig00001129
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c42 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a01,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001128
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c41 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a02,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001127
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c40 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a03,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001126
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a04,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001125
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a05,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001124
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a06,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001123
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a07,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001122
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a08,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001121
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c3a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a09,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001120
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c39 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ca,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009aa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c38 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009eb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ab,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c37 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ac,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c36 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ad,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c35 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ce,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ae,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c34 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009af,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig0000111a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c33 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig00001119
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c32 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001128,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000950
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c31 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001127,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000951
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c30 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001126,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000952
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001125,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000953
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001124,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000954
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001123,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000955
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001122,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000956
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001121,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000957
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c2a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001120,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000958
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c29 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000959
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c28 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c27 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c26 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c25 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c24 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000111a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c23 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001119,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000095f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c22 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a01,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001118
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c21 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a02,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001117
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c20 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a03,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001116
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a04,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001115
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a05,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001114
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a06,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001113
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a07,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001112
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a08,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001111
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c1a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a09,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001110
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c19 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ca,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009aa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c18 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009eb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ab,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c17 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ac,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c16 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ad,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c15 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ce,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ae,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c14 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009af,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig0000110a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c13 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig00001109
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c12 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001118,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000960
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c11 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001117,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000961
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c10 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001116,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000962
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001115,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000963
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001114,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000964
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001113,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000965
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001112,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000966
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001111,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000967
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c0a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001110,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000968
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c09 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000969
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c08 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c07 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c06 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c05 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c04 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000110a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c03 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001109,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000096f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c02 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a01,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001108
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c01 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a02,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001107
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c00 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a03,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001106
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a04,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001105
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bfe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a05,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001104
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bfd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a06,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001103
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bfc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a07,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001102
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bfb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a08,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001101
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bfa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a09,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig00001100
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ca,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009aa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009eb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ab,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ac,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ad,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010fc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ce,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ae,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010fb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009af,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001108,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000970
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001107,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000971
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bf0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001106,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000972
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001105,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000973
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001104,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000974
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001103,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000975
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001102,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000976
    );
  blk00000001_blk000001a2_blk000001a3_blk00000beb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001101,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000977
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001100,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000978
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ff,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000979
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010fe,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010fd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010fc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010fb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010fa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000097f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a01,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a02,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000be0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a03,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bdf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a04,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bde : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a05,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bdd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a06,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bdc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a07,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bdb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a08,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bda : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a09,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ca,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009aa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009eb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ab,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ac,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ad,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ce,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009ae,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a0f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009ef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009cf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009af,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a10,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009f0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009d0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009b0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010e9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000980
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000981
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bd0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000982
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bcf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000983
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000984
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bcd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000985
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bcc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000986
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bcb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000987
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010f0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000988
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ef,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000989
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ee,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ed,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ec,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010eb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ea,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010e9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000098f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010df,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010db,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bc0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010dd,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bbf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d9,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bbe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010de,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bbd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010da,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bbc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010dc,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bbb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010e0,
      Q => blk00000001_blk000001a2_blk000001a3_sig000010e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bba : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000991,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000992,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000993,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000994,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000995,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000996,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000997,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000998,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000999,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bb0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000baf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010cd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bae : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010cc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bad : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009de,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009be,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bac : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009ff,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009df,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000bab : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e3,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e4,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000baa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000910
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000911
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000912
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000913
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000914
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000915
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000916
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000917
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010d0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000918
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010cf,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000919
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ba0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ce,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010cd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010cc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010cb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ca,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000091f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b9a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000991,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b99 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000992,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b98 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000993,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b97 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000994,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b96 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000995,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b95 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000996,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b94 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000997,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b93 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000998,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b92 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000999,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b91 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b90 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010be
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009de,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009be,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009ff,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009df,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e5,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e6,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b8a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000920
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b89 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000921
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b88 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000922
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b87 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000923
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b86 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000924
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b85 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000925
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b84 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000926
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b83 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000927
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b82 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010c0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000928
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b81 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010bf,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000929
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b80 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010be,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010bd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010bc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010bb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ba,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000092f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b7a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000991,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b79 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000992,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b78 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000993,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b77 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000994,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b76 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000995,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b75 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000996,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b74 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000997,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b73 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000998,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b72 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000999,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b71 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b70 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009de,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009be,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009ff,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009df,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e7,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e8,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b6a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000930
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b69 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000931
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b68 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000932
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b67 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000933
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b66 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000934
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b65 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000935
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b64 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000936
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b63 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000937
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b62 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010b0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000938
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b61 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010af,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000939
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b60 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ae,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ad,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ac,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010ab,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010aa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000093f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b5a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000991,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b59 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000992,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b58 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000993,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b57 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000994,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b56 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000995,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b55 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000996,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b54 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000997,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b53 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000998,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b52 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009f9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009d9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009b9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000999,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig000010a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b51 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009da,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009ba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b50 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009db,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009dd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009fe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009de,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009be,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000009ff,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009df,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009bf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000099f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig0000109a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000a00,
      I1 => blk00000001_blk000001a2_blk000001a3_sig000009e0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig000009c0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig000009a0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000010e1,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000010e2,
      O => blk00000001_blk000001a2_blk000001a3_sig00001099
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b4a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000940
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b49 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000941
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b48 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000942
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b47 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000943
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b46 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000944
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b45 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000945
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b44 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000946
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b43 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000947
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b42 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000010a0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000948
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b41 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000949
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b40 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig0000109a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001099,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000094f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000b3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00001098,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000990
    );
  blk00000001_blk000001a2_blk000001a3_blk00000581 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000007f7,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000580 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c41
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c40
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000057a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fc0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000579 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fbf,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000578 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fbe,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000577 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fbd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000099a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000576 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fbc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000999
    );
  blk00000001_blk000001a2_blk000001a3_blk00000575 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fbb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000998
    );
  blk00000001_blk000001a2_blk000001a3_blk00000574 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fba,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000997
    );
  blk00000001_blk000001a2_blk000001a3_blk00000573 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000996
    );
  blk00000001_blk000001a2_blk000001a3_blk00000572 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000995
    );
  blk00000001_blk000001a2_blk000001a3_blk00000571 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000994
    );
  blk00000001_blk000001a2_blk000001a3_blk00000570 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000993
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000992
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000991
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000056d_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000056c_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000056b_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000056a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fb0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000056a_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000569 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000faf,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000569_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000568 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fae,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000568_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000567 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000566 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000565 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000564 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000563 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000562 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000561 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fc0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000560 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fbf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fbe
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fbd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b9a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fbc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b99,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b9a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fbb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b98,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b99,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b9a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fba
    );
  blk00000001_blk000001a2_blk000001a3_blk0000055a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b97,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b98,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b99,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b9a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000559 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b96,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b97,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b98,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b99,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000558 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b95,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b96,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b97,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b98,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000557 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b94,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b95,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b96,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b97,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000556 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b93,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b94,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b95,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b96,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000555 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b92,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b93,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b94,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b95,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000554 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b91,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b92,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b93,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b94,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000553 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b90,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b91,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b92,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b93,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000552 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b90,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b91,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b92,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000551 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b8f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b90,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b91,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fb0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000550 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000b8f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b90,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000faf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000b8f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fae
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fad,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c44
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fac,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c43
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fab,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c42
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000faa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000054a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000549 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000548 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000547 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000546 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000545 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000544 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000543 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000542 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000541 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000fa0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000540 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009a1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f9a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000053b_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000053a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f99,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000053a_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000539 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f98,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000539_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000538 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f97,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000538_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000537 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f96,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000537_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000536 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f95,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000536_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000535 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000534 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000533 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000532 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bba,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000faa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000531 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000530 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bb0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000052a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000baf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bb0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000529 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bae,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000baf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bb0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000528 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bad,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bae,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000baf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bb0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000fa0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000527 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bac,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bad,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bae,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000baf,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000526 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bab,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bac,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bad,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bae,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000525 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000baa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bab,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bac,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bad,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000524 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000baa,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bab,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bac,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000523 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000baa,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bab,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000522 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000baa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f9a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000521 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f99
    );
  blk00000001_blk000001a2_blk000001a3_blk00000520 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ba5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f98
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ba5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f97
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000ba5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f96
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000ba5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f95
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f94,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c47
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f93,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c46
    );
  blk00000001_blk000001a2_blk000001a3_blk0000051a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f92,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c45
    );
  blk00000001_blk000001a2_blk000001a3_blk00000519 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f91,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000518 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f90,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000517 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009be
    );
  blk00000001_blk000001a2_blk000001a3_blk00000516 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000515 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000514 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000513 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000512 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f8a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000511 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f89,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000510 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f88,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f87,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f86,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f85,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f84,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f83,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000050a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f82,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000509 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f81,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000509_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000508 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f80,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000508_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000507 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000507_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000506 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000506_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000505 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000505_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000504 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000504_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000503 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f94
    );
  blk00000001_blk000001a2_blk000001a3_blk00000502 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bfb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f93
    );
  blk00000001_blk000001a2_blk000001a3_blk00000501 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bfa,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f92
    );
  blk00000001_blk000001a2_blk000001a3_blk00000500 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfa,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f91
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfa,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f90
    );
  blk00000001_blk000001a2_blk000001a3_blk000004fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfa,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8f
    );
  blk00000001_blk000001a2_blk000001a3_blk000004fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8e
    );
  blk00000001_blk000001a2_blk000001a3_blk000004fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8d
    );
  blk00000001_blk000001a2_blk000001a3_blk000004fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8c
    );
  blk00000001_blk000001a2_blk000001a3_blk000004fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8b
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f8a
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f89
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bf0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f88
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bef,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bf0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f87
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bef,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bf0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f86
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bed,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bef,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bf0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f85
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bec,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bed,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bee,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bef,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f84
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000beb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bed,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bee,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f83
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bea,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000beb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bec,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bed,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f82
    );
  blk00000001_blk000001a2_blk000001a3_blk000004f0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000beb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bec,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f81
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ef : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bea,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000beb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f80
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ee : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bea,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7f
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ed : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7e
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ec : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7d
    );
  blk00000001_blk000001a2_blk000001a3_blk000004eb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7c
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4a
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f7a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c49
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f79,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c48
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f78,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d0
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f77,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009cf
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f76,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ce
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f75,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009cd
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f74,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009cc
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f73,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009cb
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f72,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ca
    );
  blk00000001_blk000001a2_blk000001a3_blk000004e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f71,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c9
    );
  blk00000001_blk000001a2_blk000001a3_blk000004df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f70,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c8
    );
  blk00000001_blk000001a2_blk000001a3_blk000004de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c7
    );
  blk00000001_blk000001a2_blk000001a3_blk000004dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c6
    );
  blk00000001_blk000001a2_blk000001a3_blk000004dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c5
    );
  blk00000001_blk000001a2_blk000001a3_blk000004db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c4
    );
  blk00000001_blk000001a2_blk000001a3_blk000004da : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c3
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f6a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c2
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f69,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009c1
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f68,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d7_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f67,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d6_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f66,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d5_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f65,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d4_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f64,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d3_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f63,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004d2_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7b
    );
  blk00000001_blk000001a2_blk000001a3_blk000004d0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c11,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f7a
    );
  blk00000001_blk000001a2_blk000001a3_blk000004cf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c10,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c11,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f79
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ce : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c10,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c11,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c12,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f78
    );
  blk00000001_blk000001a2_blk000001a3_blk000004cd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c10,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c11,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f77
    );
  blk00000001_blk000001a2_blk000001a3_blk000004cc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c10,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f76
    );
  blk00000001_blk000001a2_blk000001a3_blk000004cb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f75
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ca : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f74
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c0a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f73
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c09,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c0a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f72
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c08,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c09,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c0a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f71
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c07,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c08,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c09,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c0a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f70
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c06,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c07,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c08,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c09,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6f
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c05,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c06,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c07,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c08,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6e
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c04,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c05,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c06,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c07,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6d
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c03,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c04,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c05,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c06,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6c
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c02,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c03,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c04,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c05,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6b
    );
  blk00000001_blk000001a2_blk000001a3_blk000004c0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c01,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c02,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c03,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c04,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f6a
    );
  blk00000001_blk000001a2_blk000001a3_blk000004bf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c00,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c01,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c02,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c03,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f69
    );
  blk00000001_blk000001a2_blk000001a3_blk000004be : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bff,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c00,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c01,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c02,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f68
    );
  blk00000001_blk000001a2_blk000001a3_blk000004bd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bfe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bff,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c00,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c01,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f67
    );
  blk00000001_blk000001a2_blk000001a3_blk000004bc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bfd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfe,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bff,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c00,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f66
    );
  blk00000001_blk000001a2_blk000001a3_blk000004bb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bfd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfe,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bff,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f65
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ba : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bfd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfe,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f64
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bfd,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f63
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f62,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4d
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f61,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4c
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f60,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4b
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e0
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009df
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009de
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009dd
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009dc
    );
  blk00000001_blk000001a2_blk000001a3_blk000004b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f5a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009db
    );
  blk00000001_blk000001a2_blk000001a3_blk000004af : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f59,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009da
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f58,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d9
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f57,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d8
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f56,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d7
    );
  blk00000001_blk000001a2_blk000001a3_blk000004ab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f55,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d6
    );
  blk00000001_blk000001a2_blk000001a3_blk000004aa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f54,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d5
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f53,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d4
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f52,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d3
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f51,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d2
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f50,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009d1
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a5_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a4_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a3_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a2_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a1_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk000004a0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f4a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk000004a0_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f62
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bcf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f61
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bce,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bcf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f60
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bcd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bce,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bcf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bcc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bcd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bce,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bcf,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000049a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bcb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bcc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bcd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bce,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000499 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bca,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bcb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bcc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bcd,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000498 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bca,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bcb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bcc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000497 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bca,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bcb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f5a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000496 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bca,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f59
    );
  blk00000001_blk000001a2_blk000001a3_blk00000495 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f58
    );
  blk00000001_blk000001a2_blk000001a3_blk00000494 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000493 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f56
    );
  blk00000001_blk000001a2_blk000001a3_blk00000492 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f55
    );
  blk00000001_blk000001a2_blk000001a3_blk00000491 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f54
    );
  blk00000001_blk000001a2_blk000001a3_blk00000490 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f53
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bc0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f52
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bbf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bc0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f51
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bbe,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bbf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bc0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f50
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bbd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bbe,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bbf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bc0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bbc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bbd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bbe,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bbf,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000048a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bbb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bbc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bbd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bbe,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000489 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bbb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bbc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bbd,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000488 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bbb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bbc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000487 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bbb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000486 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f49,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c50
    );
  blk00000001_blk000001a2_blk000001a3_blk00000485 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f48,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000484 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f47,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c4e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000483 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f46,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000482 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f45,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000481 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f44,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000480 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f43,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ed
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f42,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ec
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f41,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009eb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f40,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ea
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000047a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000479 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000478 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000477 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f3a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000476 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f39,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000475 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f38,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000474 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f37,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000473 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f36,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000473_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000472 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f35,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000472_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000471 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f34,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000471_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000470 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f33,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000470_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f32,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000046f_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f31,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000046e_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f49
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f48
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f47
    );
  blk00000001_blk000001a2_blk000001a3_blk0000046a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f46
    );
  blk00000001_blk000001a2_blk000001a3_blk00000469 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f45
    );
  blk00000001_blk000001a2_blk000001a3_blk00000468 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f44
    );
  blk00000001_blk000001a2_blk000001a3_blk00000467 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000be0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f43
    );
  blk00000001_blk000001a2_blk000001a3_blk00000466 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bdf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000be0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f42
    );
  blk00000001_blk000001a2_blk000001a3_blk00000465 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bdf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000be0,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f41
    );
  blk00000001_blk000001a2_blk000001a3_blk00000464 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bdd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bde,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bdf,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000be0,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f40
    );
  blk00000001_blk000001a2_blk000001a3_blk00000463 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bdc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bdd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bde,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bdf,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000462 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bdb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bdc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bdd,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bde,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000461 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bda,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bdb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bdc,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bdd,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000460 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bda,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bdb,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bdc,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bda,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bdb,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd9,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bda,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f3a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd8,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd9,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f39
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd7,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd8,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f38
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd6,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd7,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f37
    );
  blk00000001_blk000001a2_blk000001a3_blk0000045a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd5,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd6,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f36
    );
  blk00000001_blk000001a2_blk000001a3_blk00000459 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd4,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd5,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f35
    );
  blk00000001_blk000001a2_blk000001a3_blk00000458 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000bd1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd3,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd4,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f34
    );
  blk00000001_blk000001a2_blk000001a3_blk00000457 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000bd1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd2,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd3,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000456 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000bd1,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd2,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000455 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000bd1,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000454 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f30,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c53
    );
  blk00000001_blk000001a2_blk000001a3_blk00000453 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c52
    );
  blk00000001_blk000001a2_blk000001a3_blk00000452 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c51
    );
  blk00000001_blk000001a2_blk000001a3_blk00000451 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a00
    );
  blk00000001_blk000001a2_blk000001a3_blk00000450 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009ff
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009fe
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f2a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009fd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f29,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009fc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f28,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009fb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f27,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009fa
    );
  blk00000001_blk000001a2_blk000001a3_blk0000044a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f26,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000449 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f25,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000448 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f24,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000447 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f23,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000446 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f22,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000445 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f21,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000444 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f20,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000443 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000442 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig000009f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000441 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000441_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000440 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000440_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000043f_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f1a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000043e_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f19,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000043d_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f18,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000043c_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f30
    );
  blk00000001_blk000001a2_blk000001a3_blk0000043a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c27,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000439 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c26,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c27,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000438 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c25,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c26,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c27,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c28,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000437 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c24,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c25,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c26,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c27,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000436 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c23,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c24,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c25,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c26,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000435 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c22,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c23,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c24,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c25,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000434 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c21,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c22,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c23,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c24,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000433 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c20,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c21,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c22,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c23,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f28
    );
  blk00000001_blk000001a2_blk000001a3_blk00000432 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c20,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c21,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c22,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000431 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c20,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c21,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000430 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c20,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f25
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f24
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f23
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c1a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f22
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c19,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c1a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f21
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c18,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c19,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c1a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f20
    );
  blk00000001_blk000001a2_blk000001a3_blk0000042a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c17,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c18,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c19,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c1a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000429 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c16,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c17,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c18,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c19,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000428 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c15,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c16,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c17,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c18,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000427 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c14,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c15,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c16,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c17,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000426 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c13,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c14,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c15,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c16,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000425 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c13,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c14,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c15,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f1a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000424 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c13,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c14,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f19
    );
  blk00000001_blk000001a2_blk000001a3_blk00000423 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c13,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f18
    );
  blk00000001_blk000001a2_blk000001a3_blk00000422 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f17,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c56
    );
  blk00000001_blk000001a2_blk000001a3_blk00000421 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f16,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c55
    );
  blk00000001_blk000001a2_blk000001a3_blk00000420 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f15,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c54
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f14,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a10
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f13,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f12,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f11,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f10,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000041a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000419 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a0a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000418 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a09
    );
  blk00000001_blk000001a2_blk000001a3_blk00000417 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a08
    );
  blk00000001_blk000001a2_blk000001a3_blk00000416 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a07
    );
  blk00000001_blk000001a2_blk000001a3_blk00000415 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f0a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a06
    );
  blk00000001_blk000001a2_blk000001a3_blk00000414 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f09,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a05
    );
  blk00000001_blk000001a2_blk000001a3_blk00000413 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f08,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a04
    );
  blk00000001_blk000001a2_blk000001a3_blk00000412 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f07,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a03
    );
  blk00000001_blk000001a2_blk000001a3_blk00000411 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f06,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a02
    );
  blk00000001_blk000001a2_blk000001a3_blk00000410 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f05,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a01
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f04,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040f_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f03,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040e_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f02,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040d_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f01,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040c_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000f00,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040b_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk0000040a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000eff,
      R => blk00000001_blk000001a2_sig00000592,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk0000040a_Q_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000409 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f17
    );
  blk00000001_blk000001a2_blk000001a3_blk00000408 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c3d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f16
    );
  blk00000001_blk000001a2_blk000001a3_blk00000407 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c3c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f15
    );
  blk00000001_blk000001a2_blk000001a3_blk00000406 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c3b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f14
    );
  blk00000001_blk000001a2_blk000001a3_blk00000405 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c3a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f13
    );
  blk00000001_blk000001a2_blk000001a3_blk00000404 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c39,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f12
    );
  blk00000001_blk000001a2_blk000001a3_blk00000403 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c38,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c3a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f11
    );
  blk00000001_blk000001a2_blk000001a3_blk00000402 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c37,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c39,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c3a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f10
    );
  blk00000001_blk000001a2_blk000001a3_blk00000401 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c36,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c38,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c39,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000400 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c35,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c36,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c37,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c38,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0e
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c34,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c35,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c36,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c37,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0d
    );
  blk00000001_blk000001a2_blk000001a3_blk000003fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c33,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c34,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c35,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c36,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0c
    );
  blk00000001_blk000001a2_blk000001a3_blk000003fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c32,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c33,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c34,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c35,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0b
    );
  blk00000001_blk000001a2_blk000001a3_blk000003fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c31,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c32,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c33,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c34,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f0a
    );
  blk00000001_blk000001a2_blk000001a3_blk000003fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c30,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c31,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c32,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c33,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f09
    );
  blk00000001_blk000001a2_blk000001a3_blk000003fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c30,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c31,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c32,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f08
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c30,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c31,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f07
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c30,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f06
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f05
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f04
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c2a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f03
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000c29,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c2a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f02
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000c29,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c2a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f01
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000c29,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c2a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000f00
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_sig00000592,
      I1 => blk00000001_blk000001a2_sig00000592,
      I2 => blk00000001_blk000001a2_sig00000592,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000c29,
      I4 => blk00000001_blk000001a2_blk000001a3_sig0000090e,
      I5 => blk00000001_blk000001a2_blk000001a3_sig0000090f,
      O => blk00000001_blk000001a2_blk000001a3_sig00000eff
    );
  blk00000001_blk000001a2_blk000001a3_blk000003f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000e28,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000efe
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000809,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e9b
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000e9b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d40
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig000011b4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e28
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000802,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000efd
    );
  blk00000001_blk000001a2_blk000001a3_blk000003eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000efd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e27
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d0e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cdf
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d0d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce0
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d0c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce1
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d0b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce2
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d0a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce3
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d09,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce4
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d08,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce5
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d07,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce6
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d06,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce7
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d05,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce8
    );
  blk00000001_blk000001a2_blk000001a3_blk000003e0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d04,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ce9
    );
  blk00000001_blk000001a2_blk000001a3_blk000003df : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d03,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cea
    );
  blk00000001_blk000001a2_blk000001a3_blk000003de : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d02,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ceb
    );
  blk00000001_blk000001a2_blk000001a3_blk000003dd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d01,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cec
    );
  blk00000001_blk000001a2_blk000001a3_blk000003dc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000d00,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ced
    );
  blk00000001_blk000001a2_blk000001a3_blk000003db : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cff,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cee
    );
  blk00000001_blk000001a2_blk000001a3_blk000003da : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a21,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d0e
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a22,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d0d
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a23,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d0c
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a24,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d0b
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a25,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d0a
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a26,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d09
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a27,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d08
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a28,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d07
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a29,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d06
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d05
    );
  blk00000001_blk000001a2_blk000001a3_blk000003d0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d04
    );
  blk00000001_blk000001a2_blk000001a3_blk000003cf : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d03
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ce : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d02
    );
  blk00000001_blk000001a2_blk000001a3_blk000003cd : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d01
    );
  blk00000001_blk000001a2_blk000001a3_blk000003cc : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a2f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d00
    );
  blk00000001_blk000001a2_blk000001a3_blk000003cb : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a30,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cff
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cfe,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ccf
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cfd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd0
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cfc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd1
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cfb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd2
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cfa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd3
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd4
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd5
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd6
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf6,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd7
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf5,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd8
    );
  blk00000001_blk000001a2_blk000001a3_blk000003c0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf4,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cd9
    );
  blk00000001_blk000001a2_blk000001a3_blk000003bf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf3,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cda
    );
  blk00000001_blk000001a2_blk000001a3_blk000003be : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf2,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cdb
    );
  blk00000001_blk000001a2_blk000001a3_blk000003bd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf1,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cdc
    );
  blk00000001_blk000001a2_blk000001a3_blk000003bc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cf0,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cdd
    );
  blk00000001_blk000001a2_blk000001a3_blk000003bb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cef,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cde
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ba : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a11,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cfe
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a12,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cfd
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a13,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cfc
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a14,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cfb
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a15,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cfa
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a16,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf9
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a17,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf8
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a18,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf7
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a19,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf6
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf5
    );
  blk00000001_blk000001a2_blk000001a3_blk000003b0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf4
    );
  blk00000001_blk000001a2_blk000001a3_blk000003af : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf3
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ae : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf2
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ad : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf1
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ac : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a1f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cf0
    );
  blk00000001_blk000001a2_blk000001a3_blk000003ab : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a20,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000cef
    );
  blk00000001_blk000001a2_blk000001a3_blk000003aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7b
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7c
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7d
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000caa,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7e
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cab,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7f
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cac,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b80
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cad,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b81
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cae,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b82
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000caf,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b83
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b84
    );
  blk00000001_blk000001a2_blk000001a3_blk000003a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b85
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b86
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b87
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b88
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b89
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000039a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000399 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000398 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cb9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000397 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cba,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000396 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000395 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b40
    );
  blk00000001_blk000001a2_blk000001a3_blk00000394 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b41
    );
  blk00000001_blk000001a2_blk000001a3_blk00000393 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b42
    );
  blk00000001_blk000001a2_blk000001a3_blk00000392 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b43
    );
  blk00000001_blk000001a2_blk000001a3_blk00000391 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c70,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b44
    );
  blk00000001_blk000001a2_blk000001a3_blk00000390 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c71,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b45
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c72,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b46
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c73,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b47
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c74,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b48
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c75,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b49
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c76,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000038a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c77,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000389 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c78,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000388 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c79,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000387 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000386 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b4f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000385 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b50
    );
  blk00000001_blk000001a2_blk000001a3_blk00000384 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b51
    );
  blk00000001_blk000001a2_blk000001a3_blk00000383 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b52
    );
  blk00000001_blk000001a2_blk000001a3_blk00000382 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c93,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b67
    );
  blk00000001_blk000001a2_blk000001a3_blk00000381 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c94,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b68
    );
  blk00000001_blk000001a2_blk000001a3_blk00000380 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c95,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b69
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c96,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c97,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c98,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c99,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000037a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b6f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000379 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b70
    );
  blk00000001_blk000001a2_blk000001a3_blk00000378 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b71
    );
  blk00000001_blk000001a2_blk000001a3_blk00000377 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b72
    );
  blk00000001_blk000001a2_blk000001a3_blk00000376 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c9f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b73
    );
  blk00000001_blk000001a2_blk000001a3_blk00000375 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b74
    );
  blk00000001_blk000001a2_blk000001a3_blk00000374 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b75
    );
  blk00000001_blk000001a2_blk000001a3_blk00000373 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b76
    );
  blk00000001_blk000001a2_blk000001a3_blk00000372 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b77
    );
  blk00000001_blk000001a2_blk000001a3_blk00000371 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b78
    );
  blk00000001_blk000001a2_blk000001a3_blk00000370 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b79
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ca6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b7a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c7f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b53
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c80,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b54
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c81,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b55
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c82,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b56
    );
  blk00000001_blk000001a2_blk000001a3_blk0000036a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c83,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000369 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c84,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b58
    );
  blk00000001_blk000001a2_blk000001a3_blk00000368 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c85,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b59
    );
  blk00000001_blk000001a2_blk000001a3_blk00000367 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c86,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000366 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c87,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000365 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c88,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000364 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c89,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000363 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000362 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b5f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000361 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b60
    );
  blk00000001_blk000001a2_blk000001a3_blk00000360 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b61
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b62
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c8f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b63
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c90,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b64
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c91,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b65
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c92,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b66
    );
  blk00000001_blk000001a2_blk000001a3_blk0000035a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c57,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000359 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c58,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000358 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c59,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000356 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000355 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000354 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000353 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000352 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c5f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000351 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c60,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b34
    );
  blk00000001_blk000001a2_blk000001a3_blk00000350 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c61,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b35
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c62,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b36
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c63,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b37
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c64,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b38
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c65,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b39
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c66,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000034a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c67,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000349 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c68,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000348 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c69,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000347 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000c6a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000346 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cbb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b17
    );
  blk00000001_blk000001a2_blk000001a3_blk00000345 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cbc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b18
    );
  blk00000001_blk000001a2_blk000001a3_blk00000344 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cbd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b19
    );
  blk00000001_blk000001a2_blk000001a3_blk00000343 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cbe,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000342 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cbf,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000341 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000340 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b1f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b20
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b21
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b22
    );
  blk00000001_blk000001a2_blk000001a3_blk0000033a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b23
    );
  blk00000001_blk000001a2_blk000001a3_blk00000339 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b24
    );
  blk00000001_blk000001a2_blk000001a3_blk00000338 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cc9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b25
    );
  blk00000001_blk000001a2_blk000001a3_blk00000337 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cca,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000336 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ccb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000335 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ccc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b28
    );
  blk00000001_blk000001a2_blk000001a3_blk00000334 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ccd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000333 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000cce,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000332 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b16,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000331 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b15,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000330 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b14,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000a9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b13,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000aa
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b12,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000ab
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b11,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000ac
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b10,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000ad
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000ae
    );
  blk00000001_blk000001a2_blk000001a3_blk0000032a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000329 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000328 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000327 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000326 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b0a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000325 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b09,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000324 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b08,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000323 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b07,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000322 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000829,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000849,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000869,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000889,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b16
    );
  blk00000001_blk000001a2_blk000001a3_blk00000321 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000828,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000848,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000868,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000888,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b15
    );
  blk00000001_blk000001a2_blk000001a3_blk00000320 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000827,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000847,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000867,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000887,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b14
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000826,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000846,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000866,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000886,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b13
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000825,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000845,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000865,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000885,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b12
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000824,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000844,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000864,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000884,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b11
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000823,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000843,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000863,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000883,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b10
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000822,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000842,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000862,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000882,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000031a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000821,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000841,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000861,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000881,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000319 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000820,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000840,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000860,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000880,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000318 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000317 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000316 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b0a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000315 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b09
    );
  blk00000001_blk000001a2_blk000001a3_blk00000314 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b08
    );
  blk00000001_blk000001a2_blk000001a3_blk00000313 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b07
    );
  blk00000001_blk000001a2_blk000001a3_blk00000312 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b06,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000311 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b05,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000310 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b04,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000b9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b03,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000ba
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b02,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000bb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b01,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000bc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000b00,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000bd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aff,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000be
    );
  blk00000001_blk000001a2_blk000001a3_blk0000030a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000afe,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000309 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000afd,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000308 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000afc,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000307 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000afb,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000306 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000afa,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000305 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af9,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000304 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af8,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000303 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af7,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_sig000000c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000302 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000819,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000839,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000859,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000879,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b06
    );
  blk00000001_blk000001a2_blk000001a3_blk00000301 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000818,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000838,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000858,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000878,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b05
    );
  blk00000001_blk000001a2_blk000001a3_blk00000300 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000817,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000837,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000857,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000877,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b04
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000816,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000836,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000856,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000876,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b03
    );
  blk00000001_blk000001a2_blk000001a3_blk000002fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000815,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000835,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000855,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000875,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b02
    );
  blk00000001_blk000001a2_blk000001a3_blk000002fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000814,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000834,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000854,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000874,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b01
    );
  blk00000001_blk000001a2_blk000001a3_blk000002fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000813,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000833,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000853,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000873,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000b00
    );
  blk00000001_blk000001a2_blk000001a3_blk000002fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000812,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000832,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000852,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000872,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aff
    );
  blk00000001_blk000001a2_blk000001a3_blk000002fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000811,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000831,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000851,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000871,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000afe
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000810,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000830,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000850,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000870,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000afd
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000afc
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000afb
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000afa
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af9
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af8
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007ec,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007eb,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af7
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a20
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1f
    );
  blk00000001_blk000001a2_blk000001a3_blk000002f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1e
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1d
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1c
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1b
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000af0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a1a
    );
  blk00000001_blk000001a2_blk000001a3_blk000002eb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aef,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a19
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aee,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a18
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aed,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a17
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aec,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a16
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aeb,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a15
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aea,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a14
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae9,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a13
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae8,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a12
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae7,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a11
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000819,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000839,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000859,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000879,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af6
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000818,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000838,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000858,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000878,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af5
    );
  blk00000001_blk000001a2_blk000001a3_blk000002e0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000817,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000837,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000857,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000877,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af4
    );
  blk00000001_blk000001a2_blk000001a3_blk000002df : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000816,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000836,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000856,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000876,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af3
    );
  blk00000001_blk000001a2_blk000001a3_blk000002de : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000815,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000835,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000855,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000875,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af2
    );
  blk00000001_blk000001a2_blk000001a3_blk000002dd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000814,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000834,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000854,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000874,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af1
    );
  blk00000001_blk000001a2_blk000001a3_blk000002dc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000813,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000833,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000853,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000873,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000af0
    );
  blk00000001_blk000001a2_blk000001a3_blk000002db : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000812,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000832,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000852,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000872,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aef
    );
  blk00000001_blk000001a2_blk000001a3_blk000002da : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000811,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000831,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000851,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000871,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aee
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000810,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000830,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000850,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000870,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aed
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aec
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aeb
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aea
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae9
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae8
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000080a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000082a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000084a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000086a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae7
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d50
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4f
    );
  blk00000001_blk000001a2_blk000001a3_blk000002d0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4e
    );
  blk00000001_blk000001a2_blk000001a3_blk000002cf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4d
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4c
    );
  blk00000001_blk000001a2_blk000001a3_blk000002cd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4b
    );
  blk00000001_blk000001a2_blk000001a3_blk000002cc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ae0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d4a
    );
  blk00000001_blk000001a2_blk000001a3_blk000002cb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000adf,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d49
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ade,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d48
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000add,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d47
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000adc,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d46
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000adb,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d45
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ada,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d44
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad9,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d43
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad8,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d42
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad7,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d41
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000839,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000859,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000879,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000819,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae6
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000838,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000858,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000878,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000818,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae5
    );
  blk00000001_blk000001a2_blk000001a3_blk000002c0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000837,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000857,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000877,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000817,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae4
    );
  blk00000001_blk000001a2_blk000001a3_blk000002bf : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000836,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000856,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000876,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000816,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae3
    );
  blk00000001_blk000001a2_blk000001a3_blk000002be : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000835,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000855,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000875,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000815,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae2
    );
  blk00000001_blk000001a2_blk000001a3_blk000002bd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000834,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000854,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000874,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000814,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae1
    );
  blk00000001_blk000001a2_blk000001a3_blk000002bc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000833,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000853,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000873,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000813,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ae0
    );
  blk00000001_blk000001a2_blk000001a3_blk000002bb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000832,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000852,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000872,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000812,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000adf
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ba : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000831,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000851,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000871,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000811,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ade
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000830,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000850,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000870,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000810,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000add
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000adc
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000adb
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ada
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad9
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad8
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000082a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000084a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000086a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000080a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad7
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc3
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc2
    );
  blk00000001_blk000001a2_blk000001a3_blk000002b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc1
    );
  blk00000001_blk000001a2_blk000001a3_blk000002af : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc0
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dbf
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ad : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dbe
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ac : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ad0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dbd
    );
  blk00000001_blk000001a2_blk000001a3_blk000002ab : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000acf,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dbc
    );
  blk00000001_blk000001a2_blk000001a3_blk000002aa : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ace,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dbb
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000acd,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dba
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000acc,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db9
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000acb,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db8
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aca,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db7
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac9,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db6
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac8,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db5
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac7,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000db4
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a2 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000859,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000879,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000819,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000839,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad6
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a1 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000858,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000878,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000818,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000838,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad5
    );
  blk00000001_blk000001a2_blk000001a3_blk000002a0 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000857,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000877,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000817,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000837,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000856,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000876,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000816,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000836,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000855,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000875,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000815,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000835,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000854,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000874,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000814,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000834,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000853,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000873,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000813,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000833,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ad0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000852,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000872,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000812,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000832,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000acf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000029a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000851,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000871,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000811,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000831,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ace
    );
  blk00000001_blk000001a2_blk000001a3_blk00000299 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000850,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000870,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000810,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000830,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000acd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000298 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000acc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000297 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000acb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000296 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000295 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000294 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000293 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000084a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000086a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000080a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000082a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000292 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e38
    );
  blk00000001_blk000001a2_blk000001a3_blk00000291 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e37
    );
  blk00000001_blk000001a2_blk000001a3_blk00000290 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e36
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e35
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e34
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e33
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ac0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e32
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000abf,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e31
    );
  blk00000001_blk000001a2_blk000001a3_blk0000028a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000abe,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000289 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000abd,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000288 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000abc,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000287 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000abb,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000286 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aba,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000285 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab9,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000284 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab8,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000283 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab7,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000282 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000879,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000819,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000839,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000859,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000281 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000878,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000818,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000838,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000858,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000280 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000877,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000817,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000837,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000857,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000876,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000816,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000836,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000856,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000875,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000815,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000835,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000855,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000874,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000814,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000834,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000854,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000873,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000813,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000833,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000853,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ac0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000872,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000812,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000832,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000852,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000abf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000027a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000871,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000811,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000831,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000851,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000abe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000279 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000870,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000810,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000830,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000850,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000abd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000278 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000abc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000277 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000abb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000276 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000275 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000274 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000273 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000086a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000080a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000082a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000084a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000272 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000271 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000270 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000ab0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a2a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aaf,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a29
    );
  blk00000001_blk000001a2_blk000001a3_blk0000026a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aae,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a28
    );
  blk00000001_blk000001a2_blk000001a3_blk00000269 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aad,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000268 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aac,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000267 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aab,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a25
    );
  blk00000001_blk000001a2_blk000001a3_blk00000266 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aaa,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a24
    );
  blk00000001_blk000001a2_blk000001a3_blk00000265 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa9,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a23
    );
  blk00000001_blk000001a2_blk000001a3_blk00000264 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa8,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a22
    );
  blk00000001_blk000001a2_blk000001a3_blk00000263 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa7,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a21
    );
  blk00000001_blk000001a2_blk000001a3_blk00000262 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000829,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000849,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000869,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000889,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000261 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000828,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000848,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000868,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000888,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000260 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000827,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000847,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000867,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000887,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000826,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000846,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000866,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000886,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000825,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000845,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000865,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000885,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000824,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000844,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000864,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000884,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000823,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000843,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000863,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000883,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000ab0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000822,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000842,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000862,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000882,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aaf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000025a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000821,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000841,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000861,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000881,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000259 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000820,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000840,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000860,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000880,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000258 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000257 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000256 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aaa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000255 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000254 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000253 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000081a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000083a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000085a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000087a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000252 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa6,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d60
    );
  blk00000001_blk000001a2_blk000001a3_blk00000251 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa5,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000250 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa4,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa3,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa2,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa1,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000aa0,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d5a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9f,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d59
    );
  blk00000001_blk000001a2_blk000001a3_blk0000024a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9e,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d58
    );
  blk00000001_blk000001a2_blk000001a3_blk00000249 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9d,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000248 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9c,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d56
    );
  blk00000001_blk000001a2_blk000001a3_blk00000247 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9b,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d55
    );
  blk00000001_blk000001a2_blk000001a3_blk00000246 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a9a,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d54
    );
  blk00000001_blk000001a2_blk000001a3_blk00000245 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a99,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d53
    );
  blk00000001_blk000001a2_blk000001a3_blk00000244 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a98,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d52
    );
  blk00000001_blk000001a2_blk000001a3_blk00000243 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a97,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000d51
    );
  blk00000001_blk000001a2_blk000001a3_blk00000242 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000849,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000869,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000889,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000829,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000241 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000848,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000868,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000888,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000828,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000240 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000847,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000867,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000887,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000827,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000846,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000866,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000886,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000826,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000845,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000865,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000885,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000825,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000844,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000864,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000884,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000824,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000843,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000863,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000883,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000823,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000aa0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000842,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000862,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000882,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000822,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000023a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000841,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000861,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000881,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000821,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000239 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000840,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000860,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000880,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000820,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000238 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000237 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000236 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a9a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000235 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a99
    );
  blk00000001_blk000001a2_blk000001a3_blk00000234 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a98
    );
  blk00000001_blk000001a2_blk000001a3_blk00000233 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000083a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000085a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000087a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000081a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a97
    );
  blk00000001_blk000001a2_blk000001a3_blk00000232 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a96,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000231 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a95,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000230 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a94,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a93,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dd0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a92,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dcf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a91,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dce
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a90,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dcd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8f,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dcc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000022a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8e,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dcb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000229 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8d,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000228 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8c,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000227 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8b,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000226 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a8a,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000225 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a89,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000224 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a88,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000223 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a87,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000dc4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000222 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000869,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000889,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000829,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000849,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a96
    );
  blk00000001_blk000001a2_blk000001a3_blk00000221 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000868,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000888,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000828,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000848,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a95
    );
  blk00000001_blk000001a2_blk000001a3_blk00000220 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000867,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000887,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000827,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000847,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a94
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021f : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000866,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000886,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000826,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000846,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a93
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021e : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000865,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000885,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000825,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000845,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a92
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021d : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000864,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000884,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000824,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000844,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a91
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021c : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000863,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000883,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000823,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000843,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a90
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021b : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000862,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000882,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000822,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000842,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000021a : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000861,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000881,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000821,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000841,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000219 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000860,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000880,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000820,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000840,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000218 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000217 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000216 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a8a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000215 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a89
    );
  blk00000001_blk000001a2_blk000001a3_blk00000214 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a88
    );
  blk00000001_blk000001a2_blk000001a3_blk00000213 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000085a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000087a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000081a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000083a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a87
    );
  blk00000001_blk000001a2_blk000001a3_blk00000212 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a86,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e48
    );
  blk00000001_blk000001a2_blk000001a3_blk00000211 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a85,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e47
    );
  blk00000001_blk000001a2_blk000001a3_blk00000210 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a84,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e46
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020f : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a83,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e45
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020e : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a82,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e44
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020d : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a81,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e43
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020c : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a80,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e42
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020b : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7f,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e41
    );
  blk00000001_blk000001a2_blk000001a3_blk0000020a : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7e,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e40
    );
  blk00000001_blk000001a2_blk000001a3_blk00000209 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7d,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000208 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7c,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000207 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7b,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000206 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a7a,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000205 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a79,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000204 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a78,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e3a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000203 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007f6,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a77,
      R => blk00000001_blk000001a2_blk000001a3_sig00000800,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000e39
    );
  blk00000001_blk000001a2_blk000001a3_blk00000202 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000889,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000829,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000849,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000869,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a86
    );
  blk00000001_blk000001a2_blk000001a3_blk00000201 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000888,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000828,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000848,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000868,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a85
    );
  blk00000001_blk000001a2_blk000001a3_blk00000200 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000887,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000827,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000847,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000867,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a84
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ff : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000886,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000826,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000846,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000866,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a83
    );
  blk00000001_blk000001a2_blk000001a3_blk000001fe : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000885,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000825,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000845,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000865,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a82
    );
  blk00000001_blk000001a2_blk000001a3_blk000001fd : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000884,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000824,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000844,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000864,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a81
    );
  blk00000001_blk000001a2_blk000001a3_blk000001fc : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000883,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000823,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000843,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000863,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a80
    );
  blk00000001_blk000001a2_blk000001a3_blk000001fb : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000882,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000822,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000842,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000862,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7f
    );
  blk00000001_blk000001a2_blk000001a3_blk000001fa : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000881,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000821,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000841,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000861,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7e
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f9 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000880,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000820,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00000840,
      I3 => blk00000001_blk000001a2_blk000001a3_sig00000860,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7d
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f8 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083f,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085f,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7c
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f7 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083e,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085e,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7b
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f6 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083d,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085d,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a7a
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f5 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083c,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085c,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a79
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f4 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083b,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085b,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a78
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f3 : LUT6
    generic map(
      INIT => X"FF00F0F0CCCCAAAA"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000087a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000081a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000083a,
      I3 => blk00000001_blk000001a2_blk000001a3_sig0000085a,
      I4 => blk00000001_blk000001a2_blk000001a3_sig000007e8,
      I5 => blk00000001_blk000001a2_blk000001a3_sig000007e7,
      O => blk00000001_blk000001a2_blk000001a3_sig00000a77
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a76,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a47
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a75,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a48
    );
  blk00000001_blk000001a2_blk000001a3_blk000001f0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a74,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a49
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ef : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a73,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4a
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ee : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a72,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4b
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ed : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a71,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4c
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ec : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a70,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4d
    );
  blk00000001_blk000001a2_blk000001a3_blk000001eb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4e
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ea : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a4f
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a50
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a51
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a52
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a6a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a53
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a69,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a54
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a68,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a55
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a67,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a56
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000073,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a76
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000072,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a75
    );
  blk00000001_blk000001a2_blk000001a3_blk000001e0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000071,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a74
    );
  blk00000001_blk000001a2_blk000001a3_blk000001df : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000070,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a73
    );
  blk00000001_blk000001a2_blk000001a3_blk000001de : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a72
    );
  blk00000001_blk000001a2_blk000001a3_blk000001dd : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a71
    );
  blk00000001_blk000001a2_blk000001a3_blk000001dc : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a70
    );
  blk00000001_blk000001a2_blk000001a3_blk000001db : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6f
    );
  blk00000001_blk000001a2_blk000001a3_blk000001da : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6e
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000006a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6d
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000069,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6c
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000068,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6b
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000067,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a6a
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000066,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a69
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000065,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a68
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000064,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a67
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a66,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a37
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d1 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a65,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a38
    );
  blk00000001_blk000001a2_blk000001a3_blk000001d0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a64,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a39
    );
  blk00000001_blk000001a2_blk000001a3_blk000001cf : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a63,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3a
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ce : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a62,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3b
    );
  blk00000001_blk000001a2_blk000001a3_blk000001cd : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a61,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3c
    );
  blk00000001_blk000001a2_blk000001a3_blk000001cc : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a60,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3d
    );
  blk00000001_blk000001a2_blk000001a3_blk000001cb : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5f,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3e
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ca : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5e,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a3f
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c9 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5d,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a40
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c8 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5c,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a41
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c7 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5b,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a42
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c6 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a5a,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a43
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c5 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a59,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a44
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c4 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a58,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a45
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c3 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a57,
      R => blk00000001_blk000001a2_sig00000592,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a46
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c2 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000083,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a66
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c1 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000082,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a65
    );
  blk00000001_blk000001a2_blk000001a3_blk000001c0 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000081,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a64
    );
  blk00000001_blk000001a2_blk000001a3_blk000001bf : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000080,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a63
    );
  blk00000001_blk000001a2_blk000001a3_blk000001be : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a62
    );
  blk00000001_blk000001a2_blk000001a3_blk000001bd : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a61
    );
  blk00000001_blk000001a2_blk000001a3_blk000001bc : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a60
    );
  blk00000001_blk000001a2_blk000001a3_blk000001bb : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5f
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ba : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5e
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b9 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig0000007a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5d
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b8 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000079,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5c
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b7 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000078,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5b
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b6 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000077,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a5a
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b5 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000076,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a59
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b4 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000075,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a58
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b3 : SRL16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_sig00000801,
      A1 => blk00000001_blk000001a2_sig00000592,
      A2 => blk00000001_blk000001a2_sig00000592,
      A3 => blk00000001_blk000001a2_sig00000592,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig00000074,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a57
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b2 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000089,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a31
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b1 : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000088,
      S => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a32
    );
  blk00000001_blk000001a2_blk000001a3_blk000001b0 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000087,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a33
    );
  blk00000001_blk000001a2_blk000001a3_blk000001af : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000086,
      S => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a34
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ae : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000085,
      R => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a35
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ad : FDSE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig0000090c,
      D => blk00000001_sig00000084,
      S => blk00000001_sig00000099,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000a36
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig0000090d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000809
    );
  blk00000001_blk000001a2_blk000001a3_blk000001ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a31,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000803
    );
  blk00000001_blk000001a2_blk000001a3_blk000001aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a32,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000804
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a33,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000805
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a34,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000806
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a35,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000807
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => aclk,
      CE => blk00000001_blk000001a2_blk000001a3_sig000007ff,
      D => blk00000001_blk000001a2_blk000001a3_sig00000a36,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000808
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a5 : GND
    port map (
      G => blk00000001_blk000001a2_sig00000592
    );
  blk00000001_blk000001a2_blk000001a3_blk000001a4 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_sig00000801
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d6 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b7a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001481
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d5 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b70,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001477
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d4 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001478
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d3 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001479
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d2 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d1 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005d0 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005cf : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b6a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ce : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b69,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005cd : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b7a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005cc : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b79,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005cb : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ced,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b78,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ca : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cec,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b77,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001470
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c9 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ceb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b76,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001471
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c8 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cea,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b75,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001472
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c7 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b74,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001473
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c6 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b73,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001474
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c5 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b72,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001475
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c4 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b71,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001476
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c3 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b68,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c2 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b67,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001480
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146b,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001456,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001455,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001454,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001453,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001452,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000105f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001451,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001060
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001450,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001061
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001062
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001063
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001064
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001065
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001066
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001067
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001449,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001068
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001448,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001069
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001447,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001446,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001445,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001444,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001457,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000106e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ac : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001443,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001480,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005ab : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001443,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001480,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005aa : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146c,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146a,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001469
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001469,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cdf,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001468
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001468,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce0,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001467
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001467,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce1,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001466
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001466,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce2,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001465
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001465,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce3,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001479,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001464
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001464,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce4,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001478,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001463
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001463,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce5,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001477,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001462
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001462,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce6,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001476,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001461
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk000005a0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001461,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce7,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001475,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001460
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001460,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce8,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001474,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ce9,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001473,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cea,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001472,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ceb,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001471,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cec,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001470,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000059a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ced,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000599 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001459
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000598 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001459,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      S => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001481,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001458
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000597 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001458,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001457
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000596 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146c,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001456
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000595 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001455
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000594 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001469,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001454
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000593 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001468,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001453
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000592 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001467,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001452
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000591 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001466,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000147a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001451
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000590 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001465,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001479,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001450
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001464,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001478,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001463,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001477,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001462,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001476,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001461,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001475,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001460,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001474,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk0000058a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001473,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000144a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000589 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145e,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001472,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001449
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000588 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145d,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001471,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001448
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000587 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145c,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001470,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001447
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000586 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001446
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000585 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000145a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig0000146e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001445
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000584 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001459,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001481,
      O => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001444
    );
  blk00000001_blk000001a2_blk000001a3_blk00000582_blk00000583 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000582_sig00001443
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000062b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b66,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig00001500
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000062a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f6
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000629 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f7
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000628 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f8
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000627 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b59,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f9
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000626 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b58,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fa
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000625 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b57,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fb
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000624 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ccf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b56,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fc
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000623 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b55,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fd
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000622 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b66,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ec
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000621 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b65,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ed
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000620 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b64,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ee
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061f : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b63,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ef
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061e : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b62,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f0
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061d : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cda,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b61,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f1
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061c : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b60,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f2
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f3
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000061a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f4
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000619 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b5d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f5
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000618 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b54,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fe
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000617 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b53,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ff
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000616 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ea,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001045
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000615 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001046
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000614 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001047
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000613 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001048
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000612 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001049
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000611 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104a
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000610 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d0,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104b
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cf,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104c
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ce,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104d
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cd,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104e
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cc,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000104f
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001050
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk0000060a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ca,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001051
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000609 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001052
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000608 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001053
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000607 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001054
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000606 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001055
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000605 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001056
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000604 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001057
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000603 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001058
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000602 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001059
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000601 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c2,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ff,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014eb
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk00000600 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c2,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ff,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ea
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ff : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014eb,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fe,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e9
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005fe : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e9,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fd,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e8
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005fd : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e8,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000ccf,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fc,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e7
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005fc : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e7,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd0,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fb,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e6
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005fb : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e6,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd1,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fa,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e5
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005fa : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e5,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd2,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f9,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e4
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e4,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd3,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f8,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e3
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e3,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd4,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f7,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e2
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e2,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd5,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f6,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e1
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e1,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd6,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f5,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e0
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd7,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f4,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014df
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014df,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd8,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f3,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014de
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014de,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cd9,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f2,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dd
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cda,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f1,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dc
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cdb,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f0,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014db
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005f0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014db,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cdc,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ef,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014da
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ef : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014da,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cdd,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ee,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d9
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ee : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ed,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d8
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ed : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d8,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      S => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig00001500,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d7
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ec : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d7,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ec,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d6
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005eb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014eb,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fe,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d5
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005ea : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e9,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fd,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d4
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e8,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fc,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d3
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e7,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fb,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d2
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e6,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014fa,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d1
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e5,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f9,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d0
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e4,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f8,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cf
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e3,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f7,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ce
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e2,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f6,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cd
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e1,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f5,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cc
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014e0,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f4,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014cb
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005e0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014df,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f3,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ca
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005df : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014de,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f2,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c9
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005de : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dd,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f1,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c8
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005dd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014dc,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014f0,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c7
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005dc : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014db,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ef,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c6
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005db : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014da,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ee,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c5
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005da : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d9,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014ed,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c4
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005d9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014d8,
      LI => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig00001500,
      O => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c3
    );
  blk00000001_blk000001a2_blk000001a3_blk000005d7_blk000005d8 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk000005d7_sig000014c2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000691 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000690 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001573
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068f : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001572
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068e : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001571
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001570
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068c : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068b : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000068a : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000689 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000688 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000687 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000686 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ce9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001569
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000685 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cea,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001568
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000684 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ceb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001567
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000683 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cec,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001566
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000682 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ced,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001565
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000681 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001564
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000680 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001563
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067f : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b70,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001583
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067e : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001584
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067d : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001585
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067c : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001586
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067b : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001587
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000067a : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001588
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000679 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b6a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cdf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001589
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000678 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b69,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000677 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001579
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000676 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b79,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cee,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000675 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b78,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ced,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000674 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b77,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cec,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000673 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b76,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ceb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000672 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b75,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cea,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000671 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b74,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000670 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b73,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001580
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066f : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b72,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001581
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066e : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b71,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ce6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001582
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b68,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b67,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001577,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001030
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000066a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001575,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001031
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000669 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001560,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001032
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000668 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001033
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000667 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001034
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000666 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001035
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000665 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001558,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001036
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000664 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001556,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001037
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000663 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001554,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001038
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000662 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001552,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001039
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000661 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001550,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000660 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154e,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154c,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154a,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001548,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001546,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000103f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001544,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001040
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000065a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001542,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001041
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000659 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001540,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001042
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000658 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001043
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000657 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001562,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001044
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000656 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001574,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001578
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000655 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001577
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000654 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001578,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001574,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001576
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000653 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001578,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001575
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000652 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001579,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001562
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000651 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001576,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001574,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001561
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000650 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001576,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001560
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001561,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001573,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001589,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001561,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001589,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155f,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001572,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001588,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001588,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155d,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001571,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001587,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000064a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155d,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001587,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000649 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155b,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001570,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001586,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001559
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000648 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000155b,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001586,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001558
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000647 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001559,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156f,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001585,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001557
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000646 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001559,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001585,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001556
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000645 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001557,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156e,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001584,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001555
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000644 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001557,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001584,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001554
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000643 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001555,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156d,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001583,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001553
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000642 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001555,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001583,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001552
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000641 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001553,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156c,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001582,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001551
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000640 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001553,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001582,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001550
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001551,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156b,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001581,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001551,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001581,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154f,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000156a,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001580,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001580,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154d,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001569,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000063a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154d,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000639 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154b,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001568,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001549
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000638 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000154b,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001548
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000637 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001549,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001567,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001547
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000636 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001549,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001546
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000635 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001547,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001566,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001545
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000634 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001547,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001544
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000633 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001545,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001565,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001543
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000632 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001545,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001542
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000631 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001543,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001564,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001541
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk00000630 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001543,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000157a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001540
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000062f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001541,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001563,
      S => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000062e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001541,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000158d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig0000153e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000062c_blk0000062d : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk0000062c_sig00001574
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f7 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b66,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000161a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000ccf,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001600
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f5 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd0,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f4 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd1,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f3 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd2,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f2 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd3,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f1 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd4,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006f0 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd5,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ef : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd6,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ee : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd7,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ed : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd8,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ec : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cd9,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006eb : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cda,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ea : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdb,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e9 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdc,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e8 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cdd,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e7 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e5 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd5,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001610
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e4 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd4,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001611
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e3 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd3,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001612
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e2 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b59,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd2,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001613
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e1 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b58,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd1,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001614
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006e0 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b57,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd0,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001615
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006df : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b56,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ccf,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001616
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006de : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b55,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001617
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006dd : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b66,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001606
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006dc : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b65,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cde,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001607
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006db : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b64,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cdd,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001608
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006da : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b63,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cdc,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001609
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d9 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b62,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cdb,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d8 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b61,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cda,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d7 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b60,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd9,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d6 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd8,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d5 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd7,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d4 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b5d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000cd6,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b54,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001618
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b53,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001619
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001604,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001602,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ed,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015eb,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e9,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001020
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001021
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001022
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001023
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015df,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001024
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001025
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015db,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001026
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001027
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001028
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001029
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d3,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cf,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cd,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cb,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ef,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000102f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006bc : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001601,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001619,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001605
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006bb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001619,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001604
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ba : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001605,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001601,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001618,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001603
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001605,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001618,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001602
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cc,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001606,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001603,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001601,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001617,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001603,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001617,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ee,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001600,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001616,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ee,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001616,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ec,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ff,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001615,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ec,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001615,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ea,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fe,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001614,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006b0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ea,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001614,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006af : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e8,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fd,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001613,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ae : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001613,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ad : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e6,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fc,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001612,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ac : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001612,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006ab : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e4,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fb,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001611,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006aa : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001611,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e2,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015fa,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001610,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e2,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001610,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015df
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e0,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f9,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015de
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015e0,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015de,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f8,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015de,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015db
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dc,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f7,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015da
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015dc,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015da,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f6,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk000006a0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015da,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d8,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f5,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d6,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f4,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000160a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d4,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f3,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001609,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk0000069a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001609,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000699 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d2,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f2,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001608,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000698 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d2,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001608,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000697 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d0,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f1,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001607,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000696 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015d0,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001607,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000695 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ce,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015f0,
      S => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000161a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000694 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015ce,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000692_sig0000161a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000692_sig000015cb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000692_blk00000693 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000692_sig00001601
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000074c : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001699
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000074b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b84,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b34,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168f
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000074a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b83,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b33,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001690
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000749 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b82,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b32,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001691
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000748 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b81,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b31,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001692
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000747 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b80,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b30,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001693
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000746 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001694
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000745 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001695
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000744 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001696
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000743 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001685
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000742 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001686
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000741 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001687
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000740 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001688
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073f : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001689
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073e : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b89,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b39,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168a
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073d : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b88,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b38,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168b
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073c : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b87,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b37,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168c
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b86,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b36,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168d
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000073a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b85,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b35,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168e
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000739 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001697
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000738 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b2b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001698
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000737 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001683,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff1
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000736 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff2
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000735 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff3
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000734 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff4
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000733 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff5
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000732 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff6
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000731 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001669,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff7
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000730 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001668,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff8
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001667,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff9
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001666,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ffa
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001665,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ffb
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001664,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ffc
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001663,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ffd
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000072a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001662,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ffe
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000729 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001661,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fff
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000728 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001660,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001000
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000727 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001001
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000726 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001002
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000725 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001003
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000724 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001004
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000723 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001005
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000722 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b7b,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001698,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001684
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000721 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165b,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001698,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001683
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000720 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001684,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b7c,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001697,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001682
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001682,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b7d,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001696,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001681
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001681,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b7e,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001695,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001680
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001680,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b7f,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001694,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167f
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b80,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001693,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167e
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b81,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001692,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167d
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000071a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b82,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001691,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167c
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000719 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b83,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001690,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167b
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000718 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b84,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167a
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000717 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b85,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168e,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001679
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000716 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001679,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b86,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168d,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001678
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000715 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001678,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b87,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168c,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001677
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000714 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001677,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b88,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168b,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001676
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000713 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001676,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b89,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168a,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001675
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000712 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001675,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b8a,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001689,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001674
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000711 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001674,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b8b,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001688,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001673
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000710 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001673,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b8c,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001687,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001672
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001672,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b8d,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001686,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001671
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001671,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      S => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001699,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001670
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001670,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001685,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166f
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001684,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001697,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166e
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001682,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001696,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166d
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk0000070a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001681,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001695,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166c
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000709 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001680,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001694,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166b
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000708 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167f,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001693,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000166a
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000707 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167e,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001692,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001669
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000706 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167d,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001691,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001668
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000705 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167c,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001690,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001667
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000704 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167b,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168f,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001666
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000703 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000167a,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168e,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001665
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000702 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001679,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168d,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001664
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000701 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001678,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168c,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001663
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk00000700 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001677,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168b,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001662
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006ff : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001676,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000168a,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001661
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006fe : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001675,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001689,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001660
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006fd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001674,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001688,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165f
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006fc : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001673,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001687,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165e
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006fb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001672,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001686,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165d
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006fa : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001671,
      LI => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig00001699,
      O => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165c
    );
  blk00000001_blk000001a2_blk000001a3_blk000006f8_blk000006f9 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk000006f8_sig0000165b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk000007a1 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001718
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk000007a0 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b20,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b48,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079f : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b47,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079e : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b46,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001710
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079d : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b45,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001711
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079c : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b44,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001712
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079b : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b43,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001713
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000079a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b1a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b42,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001714
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000799 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b19,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b41,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001715
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000798 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b2a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001704
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000797 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b29,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b51,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001705
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000796 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b28,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b50,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001706
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000795 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b27,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001707
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000794 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b26,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001708
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000793 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b25,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4d,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001709
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000792 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b24,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4c,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000791 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b23,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4b,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000790 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b22,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b4a,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078f : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b21,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b49,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078e : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b18,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b40,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001716
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078d : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b17,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b3f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001717
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001702,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001006
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ed,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001007
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000078a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ec,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001008
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000789 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016eb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001009
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000788 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ea,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000787 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e9,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000786 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e8,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000785 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e7,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000784 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e6,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000783 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e5,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000100f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000782 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001010
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000781 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001011
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000780 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001012
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001013
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001014
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016df,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001015
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016de,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001016
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001017
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000077a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001018
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000779 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016db,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001019
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000778 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ee,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000101a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000777 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016da,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b17,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001717,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001703
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000776 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016da,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001717,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001702
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000775 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001703,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b18,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001716,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001701
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000774 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001701,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b19,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001715,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001700
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000773 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001700,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1a,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001714,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ff
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000772 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ff,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1b,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001713,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fe
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000771 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fe,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1c,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001712,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000770 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1d,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001711,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1e,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001710,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fb,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b1f,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fa
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fa,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b20,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b21,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f8,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b22,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000076a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f7,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b23,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000769 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f6,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b24,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000768 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f5,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b25,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001709,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000767 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f4,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b26,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001708,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000766 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f3,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b27,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001707,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000765 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f2,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b28,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001706,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000764 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f1,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b29,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001705,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000763 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00000b2a,
      S => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001718,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ef
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000762 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ef,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001704,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ee
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000761 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001703,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001716,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ed
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000760 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001701,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001715,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ec
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001700,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001714,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016eb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ff,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001713,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016ea
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fe,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001712,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fd,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001711,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fc,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001710,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000075a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fb,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000759 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016fa,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000758 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f9,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000757 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f8,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000756 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f7,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000755 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f6,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig0000170a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000754 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f5,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001709,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016e0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000753 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f4,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001708,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016df
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000752 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f3,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001707,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016de
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000751 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f2,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001706,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk00000750 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f1,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001705,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016dc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000074f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016f0,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig00001718,
      O => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016db
    );
  blk00000001_blk000001a2_blk000001a3_blk0000074d_blk0000074e : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk0000074d_sig000016da
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000809 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001083,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017aa
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000808 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001791
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000807 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001790
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000806 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178f
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000805 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178e
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000804 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178d
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000803 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b80,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178c
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000802 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b81,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178b
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000801 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b82,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178a
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk00000800 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b83,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001789
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ff : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b84,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001788
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007fe : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b85,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001787
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007fd : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b86,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001786
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007fc : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b87,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001785
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007fb : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b88,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001784
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007fa : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b89,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001783
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f9 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001782
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f8 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001781
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f7 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001780
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f6 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177f
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f5 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177e
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f4 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b84,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001079,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a0
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f3 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b83,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001078,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a1
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f2 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b82,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001077,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a2
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f1 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b81,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001076,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a3
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007f0 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b80,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001075,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a4
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ef : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001074,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a5
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ee : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001073,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a6
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ed : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001072,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a7
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ec : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001083,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b8e,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001796
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007eb : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001082,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001797
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ea : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001081,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001798
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e9 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001080,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001799
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e8 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b8a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179a
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e7 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b89,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107e,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179b
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e6 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b88,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107d,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179c
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e5 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b87,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107c,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179d
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e4 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b86,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107b,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179e
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e3 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b85,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000107a,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179f
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e2 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001071,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a8
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e1 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b7b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001070,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a9
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001794,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fdc
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001792,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fdd
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fde
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001779,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fdf
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001777,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe0
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001775,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe1
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001773,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe2
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001771,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe3
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe4
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe5
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe6
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001769,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe7
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001767,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe8
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001765,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fe9
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001763,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fea
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001761,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000feb
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fec
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fed
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fee
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001759,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fef
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ff0
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007cb : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001791,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a9,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001795
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ca : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a9,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001794
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001795,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001790,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a8,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001793
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001795,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a8,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001792
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175a,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001796,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177d
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001793,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178f,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a7,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177c
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001793,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a7,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177b
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177c,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178e,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a6,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177a
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177c,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a6,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001779
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177a,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178d,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a5,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001778
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177a,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a5,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001777
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007c0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001778,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178c,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a4,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001776
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007bf : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001778,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a4,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001775
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007be : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001776,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178b,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a3,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001774
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007bd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001776,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a3,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001773
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007bc : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001774,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000178a,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a2,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001772
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007bb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001774,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a2,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001771
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ba : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001772,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001789,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a1,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001770
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001772,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a1,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176f
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001770,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001788,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a0,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176e
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001770,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017a0,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176d
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176e,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001787,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176c
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176e,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179f,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176b
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176c,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001786,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179e,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176a
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176c,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179e,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001769
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176a,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001785,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179d,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001768
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000176a,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179d,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001767
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007b0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001768,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001784,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179c,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001766
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007af : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001768,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179c,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001765
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ae : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001766,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001783,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179b,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001764
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ad : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001766,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179b,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001763
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ac : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001764,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001782,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179a,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001762
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007ab : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001764,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000179a,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001761
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007aa : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001762,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001781,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001799,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001760
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001762,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001799,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175f
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001760,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001780,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001798,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175e
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001760,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001798,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175d
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175e,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177f,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001797,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175c
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175e,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001797,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175b
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175c,
      DI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000177e,
      S => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017aa,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175a
    );
  blk00000001_blk000001a2_blk000001a3_blk000007a2_blk000007a3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig0000175c,
      LI => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig000017aa,
      O => blk00000001_blk000001a2_blk000001a3_blk000007a2_sig00001759
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000871 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001097,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000870 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001823
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086f : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b40,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001822
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086e : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b41,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001821
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b42,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001820
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086c : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b43,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086b : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b44,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000086a : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b45,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000869 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b46,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000868 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b47,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000867 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b48,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000866 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b49,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001819
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000865 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001818
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000864 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001817
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000863 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001816
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000862 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001815
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000861 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001814
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000860 : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001813
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085f : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b50,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001812
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085e : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b51,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001811
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085d : LUT2
    generic map(
      INIT => X"8"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001810
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085c : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b48,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001832
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085b : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b47,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001833
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000085a : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b46,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001834
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000859 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b45,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001835
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000858 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b44,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001089,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001836
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000857 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b43,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001088,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001837
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000856 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b42,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001087,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001838
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000855 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b41,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001086,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001839
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000854 : LUT3
    generic map(
      INIT => X"9A"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001097,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000b52,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001828
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000853 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b51,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001096,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001829
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000852 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b50,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001095,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000851 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001094,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000850 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001093,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084f : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001092,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084e : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001091,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084d : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001090,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084c : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b4a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001830
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084b : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b49,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig0000108e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001831
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000084a : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b40,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001085,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000849 : LUT3
    generic map(
      INIT => X"B4"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00000b3f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      I2 => blk00000001_blk000001a2_blk000001a3_sig00001084,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000848 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001826,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fc7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000847 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001824,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fc8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000846 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fc9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000845 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fca
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000844 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001809,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fcb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000843 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001807,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fcc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000842 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001805,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fcd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000841 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001803,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fce
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000840 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001801,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fcf
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ff,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000083a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000839 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000838 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000837 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ef,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000836 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ed,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fd9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000835 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017eb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fda
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000834 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000fdb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000833 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001823,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001827
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000832 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_sig0000106f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001826
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000831 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001827,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001822,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001825
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000830 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001827,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001824
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ec,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001828,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001825,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001821,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001839,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001825,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001839,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180e,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001820,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001838,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180e,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001838,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000082a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180c,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181f,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001837,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000829 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180c,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001837,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001809
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000828 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180a,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181e,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001836,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001808
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000827 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000180a,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001836,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001807
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000826 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001808,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181d,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001835,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001806
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000825 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001808,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001835,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001805
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000824 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001806,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181c,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001834,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001804
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000823 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001806,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001834,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001803
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000822 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001804,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181b,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001833,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001802
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000821 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001804,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001833,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001801
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000820 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001802,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000181a,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001832,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001800
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001802,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001832,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ff
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001800,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001819,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001831,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fe
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001800,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001831,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fd
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fe,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001818,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001830,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fc
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fe,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001830,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fb
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000081a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fc,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001817,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fa
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000819 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fc,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f9
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000818 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fa,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001816,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f8
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000817 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017fa,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f7
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000816 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f8,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001815,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f6
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000815 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f8,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f5
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000814 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f6,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001814,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f4
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000813 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f6,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f3
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000812 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f4,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001813,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f2
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000811 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f4,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f1
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk00000810 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f2,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001812,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f0
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000080f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f2,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000182a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ef
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000080e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f0,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001811,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001829,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ee
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000080d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017f0,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001829,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ed
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000080c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ee,
      DI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig00001810,
      S => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ec
    );
  blk00000001_blk000001a2_blk000001a3_blk0000080a_blk0000080b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017ee,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig0000183c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000080a_sig000017eb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ca : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001044,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001044,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001896
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001043,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fef,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001897
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c7 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001042,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fee,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001898
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001041,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fed,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001899
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001040,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fec,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000feb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fea,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008c0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008bf : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008be : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001039,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008bd : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001038,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008bc : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001037,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008bb : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001036,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ba : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001035,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001034,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001033,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b7 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001032,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fde,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001031,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001030,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001880,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001895,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001894,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001893,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001892,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001891,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001890,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bda
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bdb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bdc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bdd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001889,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bde
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001888,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bdf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001887,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001886,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001885,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001884,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001883,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk000008a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001882,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001881,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000187f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001030,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018aa,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bf,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001031,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018be
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018be,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001032,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001033,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000089a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001034,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000899 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bb,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001035,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000898 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ba,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001036,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000897 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001037,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000896 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b8,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001038,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000895 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b7,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001039,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000894 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000893 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000892 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000891 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b3,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000890 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b2,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b1,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001040,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018af,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001041,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001899,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ae,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001042,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001898,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ad,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001043,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001897,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000088a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ac,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001044,
      S => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018c0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000889 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bf,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001895
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000888 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018be,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001894
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000887 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bd,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001893
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000886 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bc,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001892
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000885 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018bb,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001891
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000884 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ba,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001890
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000883 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b9,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000882 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000881 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b7,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000880 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018a0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000188a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001889
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b2,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001888
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b1,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001887
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk0000087a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018b0,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000189a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001886
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000879 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018af,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001899,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001885
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000878 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ae,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001898,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001884
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000877 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ad,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001897,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001883
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000876 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ac,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018c0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001882
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000875 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018ab,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001896,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001881
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000874 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000187f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000872_sig000018aa,
      O => blk00000001_blk000001a2_blk000001a3_blk00000872_sig00001880
    );
  blk00000001_blk000001a2_blk000001a3_blk00000872_blk00000873 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000872_sig0000187f
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000923 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdb,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001944
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000922 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdb,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191a
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000921 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fda,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191b
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000920 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd9,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191c
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd8,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191d
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd7,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191e
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd6,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191f
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001029,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd5,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001920
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001028,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd4,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001921
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000091a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001027,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd3,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001922
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000919 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001026,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd2,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001923
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000918 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001025,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd1,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001924
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000917 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001024,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd0,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001925
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000916 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001023,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcf,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001926
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000915 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001022,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fce,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001927
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000914 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001021,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcd,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001928
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000913 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001020,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcc,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001929
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000912 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcb,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192a
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000911 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fca,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192b
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000910 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc9,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192c
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc8,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192d
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc7,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192e
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001904,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bbb
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001919,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bbc
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001918,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bbd
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk0000090a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001917,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bbe
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000909 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001916,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bbf
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000908 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001915,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc0
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000907 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001914,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc1
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000906 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001913,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc2
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000905 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001912,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc3
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000904 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001911,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc4
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000903 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001910,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc5
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000902 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc6
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000901 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc7
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk00000900 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc8
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bc9
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bca
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bcb
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001909,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bcc
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001908,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bcd
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001907,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bce
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001906,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bcf
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001905,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bd0
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001903,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101b,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192e,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001943
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001943,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101c,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192d,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001942
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001942,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101d,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192c,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001941
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001941,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101e,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192b,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001940
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001940,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101f,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192a,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193f
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001020,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001929,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193e
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001021,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001928,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193d
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008f0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001022,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001927,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193c
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ef : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001023,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001926,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193b
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ee : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001024,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001925,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193a
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ed : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001025,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001924,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001939
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ec : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001939,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001026,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001923,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001938
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008eb : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001938,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001027,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001922,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001937
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ea : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001937,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001028,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001921,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001936
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001936,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001029,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001920,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001935
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001935,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102a,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191f,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001934
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001934,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102b,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191e,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001933
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001933,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102c,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191d,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001932
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001932,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102d,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191c,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001931
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001931,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102e,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191b,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001930
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001930,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      S => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001944,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192f
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001943,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192d,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001919
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001942,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192c,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001918
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008e0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001941,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192b,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001917
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008df : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001940,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192a,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001916
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008de : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193f,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001929,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001915
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008dd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193e,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001928,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001914
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008dc : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193d,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001927,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001913
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008db : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193c,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001926,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001912
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008da : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193b,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001925,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001911
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000193a,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001924,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001910
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001939,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001923,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190f
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001938,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001922,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190e
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001937,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001921,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190d
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001936,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001920,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190c
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001935,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191f,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190b
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001934,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191e,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000190a
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001933,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191d,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001909
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001932,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191c,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001908
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008d0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001931,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191b,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001907
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008cf : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001930,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001944,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001906
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008ce : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192f,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000191a,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001905
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008cd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001903,
      LI => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig0000192e,
      O => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001904
    );
  blk00000001_blk000001a2_blk000001a3_blk000008cb_blk000008cc : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk000008cb_sig00001903
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000097c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000101a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000097b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000101a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000097a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001019,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000979 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001018,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000978 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001017,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000977 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001016,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000976 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001069,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001015,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000975 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001068,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001014,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000974 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001067,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001013,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000973 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001066,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001012,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000972 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001065,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001011,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000971 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001064,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001010,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000970 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001063,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096f : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001062,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096e : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001061,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096d : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001060,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096c : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096b : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000096a : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001009,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019af
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000969 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001008,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000968 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001007,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000967 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001006,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000966 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001988,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000965 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000964 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000963 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000962 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000961 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001999,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000960 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001998,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001997,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001996,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001995,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001994,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001993,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c34
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000095a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001992,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c35
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000959 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001991,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c36
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000958 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001990,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c37
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000957 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c38
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000956 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c39
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000955 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000954 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000953 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000952 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000951 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001989,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000950 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001987,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c7,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019af,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ae,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c3,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ad,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000094a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c2,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001060,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ac,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000949 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c1,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001061,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ab,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000948 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001062,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019aa,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000947 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bf,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001063,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019be
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000946 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019be,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001064,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000945 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001065,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000944 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001066,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000943 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bb,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001067,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000942 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ba,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001068,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000941 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001069,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000940 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b8,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b7,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c7,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000093a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000939 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019af,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000938 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ae,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000937 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ad,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001999
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000936 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c2,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ac,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001998
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000935 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c1,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ab,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001997
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000934 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c0,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019aa,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001996
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000933 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bf,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001995
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000932 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019be,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001994
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000931 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bd,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001993
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000930 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bc,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001992
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019bb,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001991
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019ba,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001990
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b9,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b7,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk0000092a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019a0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000929 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000928 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019c8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000198a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000927 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig0000199e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001989
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000926 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001987,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000924_sig000019b2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001988
    );
  blk00000001_blk000001a2_blk000001a3_blk00000924_blk00000925 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000924_sig00001987
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001059,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001005,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001059,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001005,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a22
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001058,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001004,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a23
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001057,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001003,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a24
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001056,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001002,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a25
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009d0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001055,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001001,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a26
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009cf : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001054,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001000,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a27
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ce : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001053,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fff,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a28
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009cd : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001052,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffe,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a29
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009cc : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001051,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffd,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009cb : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001050,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffc,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ca : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffb,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c9 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffa,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c8 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff9,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c7 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff8,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c6 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff7,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a30
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c5 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff6,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a31
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c4 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001049,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff5,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a32
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c3 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001048,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff4,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a33
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c2 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001047,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff3,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a34
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c1 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001046,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff2,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a35
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009c0 : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001045,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff1,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a36
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c13
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a21,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c14
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a20,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c15
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c16
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c17
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c18
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c19
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a19,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a18,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a17,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a16,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c1f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a15,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c20
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a14,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c21
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a13,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c22
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a12,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c23
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a11,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c24
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a10,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c25
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c26
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c27
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c28
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001045,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a36,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001046,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a35,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001047,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a34,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a49
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a49,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001048,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a33,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a48
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a48,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001049,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a32,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a47
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a47,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104a,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a31,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a46
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a46,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104b,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a30,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a45
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a45,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104c,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a44
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a44,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104d,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a43
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk000009a0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a43,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104e,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a42
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a42,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104f,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a41
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a41,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001050,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a40
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a40,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001051,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001052,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a29,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001053,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a28,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000099a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001054,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a27,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000999 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001055,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a26,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000998 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001056,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a25,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000997 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001057,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a24,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a39
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000996 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a39,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001058,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a23,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a38
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000995 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a38,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001059,
      S => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a37
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000994 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4b,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a35,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a21
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000993 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4a,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a34,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a20
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000992 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a49,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a33,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000991 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a48,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a32,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000990 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a47,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a31,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a46,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a30,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a45,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2f,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1b
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a44,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2e,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a1a
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a43,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2d,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a19
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a42,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a18
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000098a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a41,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2b,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a17
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000989 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a40,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a2a,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a16
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000988 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3f,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a29,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a15
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000987 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3e,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a28,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a14
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000986 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3d,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a27,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a13
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000985 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3c,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a26,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a12
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000984 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3b,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a25,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a11
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000983 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a3a,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a24,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a10
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000982 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a39,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a23,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0f
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000981 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a38,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a4c,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0e
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk00000980 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a37,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a22,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0d
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000097f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0b,
      LI => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a36,
      O => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0c
    );
  blk00000001_blk000001a2_blk000001a3_blk0000097d_blk0000097e : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk0000097d_sig00001a0b
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a2e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001044,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ad0
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a2d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001044,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa6
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a2c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001043,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fef,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa7
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a2b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001042,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fee,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa8
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a2a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001041,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fed,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa9
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a29 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001040,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fec,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaa
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a28 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000feb,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aab
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a27 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fea,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aac
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a26 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe9,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aad
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a25 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe8,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aae
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a24 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe7,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaf
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a23 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000103a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe6,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab0
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a22 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001039,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe5,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab1
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a21 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001038,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe4,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab2
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a20 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001037,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe3,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab3
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001036,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe2,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab4
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001035,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe1,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab5
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001034,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fe0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab6
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001033,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdf,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab7
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001032,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fde,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab8
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a1a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001031,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdd,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab9
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a19 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001030,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdc,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aba
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a18 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a8f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001030,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aba,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acf
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a17 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acf,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001031,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab9,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ace
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a16 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ace,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001032,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab8,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acd
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a15 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001033,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab7,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acc
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a14 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001034,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab6,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acb
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a13 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acb,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001035,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab5,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aca
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a12 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aca,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001036,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab4,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac9
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a11 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001037,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab3,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac8
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a10 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac8,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001038,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab2,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac7
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac7,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001039,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab1,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac6
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103a,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac5
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103b,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaf,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac4
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103c,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aae,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac3
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac3,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103d,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aad,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac2
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a0a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac2,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103e,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aac,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac1
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a09 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac1,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000103f,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aab,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac0
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a08 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001040,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaa,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abf
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a07 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abf,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001041,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa9,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abe
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a06 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abe,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001042,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa8,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abd
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a05 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001043,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa7,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abc
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a04 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001044,
      S => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ad0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abb
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a03 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acf,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab9,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa5
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a02 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ace,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab8,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa4
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a01 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acd,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab7,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa3
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk00000a00 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acc,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab6,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa2
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ff : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001acb,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab5,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa1
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009fe : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aca,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab4,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa0
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009fd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac9,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab3,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9f
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009fc : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac8,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab2,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9e
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009fb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac7,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab1,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9d
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009fa : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac6,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ab0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9c
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac5,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaf,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9b
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac4,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aae,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9a
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac3,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aad,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a99
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac2,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aac,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a98
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac1,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aab,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a97
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ac0,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aaa,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a96
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abf,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa9,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a95
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abe,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa8,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a94
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abd,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa7,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a93
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009f0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abc,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001ad0,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a92
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ef : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001abb,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa6,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a91
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ee : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a8f,
      LI => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aba,
      O => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a90
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a91,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bba
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a92,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb9
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a93,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb8
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a94,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb7
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a95,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb6
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a96,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb5
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a97,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb4
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a98,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb3
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a99,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb2
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb1
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bb0
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000baf
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bae
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bad
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a9f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bac
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bab
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000baa
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba9
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba8
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba7
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001aa5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba6
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a90,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba5
    );
  blk00000001_blk000001a2_blk000001a3_blk000009d6_blk000009d7 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk000009d6_sig00001a8f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a87 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b54
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a86 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fdb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a85 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fda,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a84 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a83 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a82 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a81 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000102a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a80 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001029,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001028,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001027,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001026,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001025,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b34
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001024,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fd0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b35
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a7a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001023,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b36
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a79 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001022,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fce,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b37
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a78 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001021,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b38
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a77 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001020,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b39
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a76 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fcb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a75 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fca,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a74 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a73 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a72 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000101b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fc7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a71 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b13,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b53
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a70 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b53,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b52
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b52,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b51
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b51,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b50
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b50,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000101f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001020,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b39,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001021,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b38,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a6a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001022,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b37,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a69 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001023,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b36,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a68 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001024,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b35,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a67 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001025,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b34,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b49
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a66 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b49,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001026,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b33,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b48
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a65 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b48,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001027,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b32,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b47
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a64 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b47,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001028,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b31,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b46
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a63 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b46,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001029,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b30,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b45
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a62 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b45,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b44
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a61 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b44,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b43
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a60 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b43,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b42
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b42,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b41
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b41,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b40
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b40,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000102f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b54,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b53,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b52,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b28
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a5a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b51,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a59 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b50,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a58 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b39,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b25
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a57 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4e,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b38,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b24
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a56 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4d,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b37,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b23
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a55 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4c,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b36,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b22
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a54 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b35,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b21
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a53 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b4a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b34,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b20
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a52 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b49,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b33,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a51 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b48,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b32,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a50 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b47,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b31,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b46,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b30,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b45,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b44,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b43,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b19
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b42,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b18
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a4a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b41,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b17
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a49 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b40,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b54,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b16
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a48 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b2a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b15
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a47 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b13,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b3e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b14
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a46 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b15,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a45 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b16,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a44 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b17,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a43 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b18,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a42 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b19,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000ba0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a41 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a40 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b1f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b9a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b20,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b99
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a3a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b21,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b98
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a39 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b22,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b97
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a38 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b23,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b96
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a37 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b24,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b95
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a36 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b25,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b94
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a35 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b26,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b93
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a34 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b27,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b92
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a33 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b28,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b91
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a32 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b29,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b90
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a31 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b14,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000b8f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a2f_blk00000a30 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000a2f_sig00001b13
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ae0 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000101a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000adf : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000101a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ade : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001019,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000add : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001018,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000adc : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001017,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000adb : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000106a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001016,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ada : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001069,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001015,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad9 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001068,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001014,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001067,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001013,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad7 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001066,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001012,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad6 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001065,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001011,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001064,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001010,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad4 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001063,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad3 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001062,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001061,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad1 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001060,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ad0 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000acf : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig0000100a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ace : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001009,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000acd : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001008,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000acc : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001007,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000acb : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000105a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001006,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aca : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b97,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd7,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbe,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd3,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000105f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac4 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd2,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001060,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac3 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd1,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001061,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd0,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001062,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bba,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcf,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001063,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bce
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ac0 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bce,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001064,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000abf : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcd,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001065,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000abe : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcc,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001066,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000abd : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcb,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001067,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000abc : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bca,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001068,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000abb : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc9,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001069,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aba : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc8,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc7,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc6,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc5,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab6 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc4,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000106e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd7,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bad
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbe,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000ab0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd2,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aaf : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd1,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bbb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aae : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd0,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bba,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aad : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcf,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aac : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bce,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aab : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcd,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aaa : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcc,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bcb,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bca,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa7 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc9,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc7,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc6,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bb0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc4,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bd8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bae,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b99
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000aa0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b97,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bc2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b98
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b99,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c12
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c11
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c10
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a9a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b9f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a98 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a97 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c0a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a96 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c09
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a95 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c08
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a94 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c07
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a93 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c06
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a92 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c05
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a91 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c04
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a90 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c03
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001ba9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c02
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001baa,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c01
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bab,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000c00
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bac,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bff
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001bad,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bfe
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a8a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b98,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bfd
    );
  blk00000001_blk000001a2_blk000001a3_blk00000a88_blk00000a89 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000a88_sig00001b97
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b39 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001059,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001005,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b38 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001059,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001005,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b37 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001058,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001004,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b36 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001057,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001003,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c34
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b35 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001056,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001002,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c35
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b34 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001055,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001001,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c36
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b33 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001054,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001000,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c37
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b32 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001053,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000fff,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c38
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b31 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001052,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffe,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c39
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b30 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001051,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001050,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104f,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104e,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ffa,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104d,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff9,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104c,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff8,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b2a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104b,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c40
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b29 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000104a,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c41
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b28 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001049,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff5,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c42
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b27 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001048,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff4,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c43
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b26 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001047,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff3,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c44
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b25 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001046,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff2,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c45
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b24 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001045,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00000ff1,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c46
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b23 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001045,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c46,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b22 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001046,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c45,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b21 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001047,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c44,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c59
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b20 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c59,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001048,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c43,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c58
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c58,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001049,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c42,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c57,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104a,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c41,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c56
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c56,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104b,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c40,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c55
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c55,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104c,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c54
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c54,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104d,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c53
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b1a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c53,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c52
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b19 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c52,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000104f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c51
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b18 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c51,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001050,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c50
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b17 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c50,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001051,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b16 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4f,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001052,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c39,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b15 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4e,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001053,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c38,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b14 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4d,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001054,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c37,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b13 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001055,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c36,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b12 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001056,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c35,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b11 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001057,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c34,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c49
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b10 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c49,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001058,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c33,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c48
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c48,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001059,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c47
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c45,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c44,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c59,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c43,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c58,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c42,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b0a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c57,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c41,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b09 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c56,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c40,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b08 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c55,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b07 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c54,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b06 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c53,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c29
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b05 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c52,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c28
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b04 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c51,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b03 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c50,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c3a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b02 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4f,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c39,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c25
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b01 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4e,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c38,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c24
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000b00 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4d,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c37,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c23
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aff : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4c,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c36,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c22
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000afe : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c35,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c21
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000afd : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c4a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c34,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c20
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000afc : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c49,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c33,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000afb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c48,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c5c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000afa : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c47,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c32,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af9 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c46,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bfc
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bfb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bfa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c20,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c21,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c22,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c23,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c24,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000af0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c25,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c26,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c27,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c28,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf1
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c29,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bf0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aeb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000aea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bec
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000beb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c2f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000bea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c30,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c31,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000be7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ae1_blk00000ae2 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ae1_sig00001c1b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c50 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c68,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000090a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c4f : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c67,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c66,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c66,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c66,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007fe,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c68,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c4f_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c4e : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c67
    );
  blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_blk00000c4d : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000c4b_blk00000c4c_sig00001c66
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000009a,
      RDCLK => aclk,
      WREN => blk00000001_sig0000009a,
      RDEN => blk00000001_sig0000009a,
      WRCLK => aclk,
      SSR => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DIP(3) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DIP(2) => blk00000001_blk000001a2_blk000001a3_sig000008a4,
      DIP(1) => blk00000001_blk000001a2_blk000001a3_sig0000089b,
      DIP(0) => blk00000001_blk000001a2_blk000001a3_sig00000892,
      DOP(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb4,
      DOP(1) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb3,
      DOP(0) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb2,
      WE(3) => blk00000001_blk000001a2_blk000001a3_sig000007ca,
      WE(2) => blk00000001_blk000001a2_blk000001a3_sig000007ca,
      WE(1) => blk00000001_blk000001a2_blk000001a3_sig000007ca,
      WE(0) => blk00000001_blk000001a2_blk000001a3_sig000007ca,
      DO(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d73_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cad,
      DO(27) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cae,
      DO(26) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caf,
      DO(25) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb0,
      DO(24) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb1,
      DO(23) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca5,
      DO(22) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca6,
      DO(21) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca7,
      DO(20) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca8,
      DO(19) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca9,
      DO(18) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caa,
      DO(17) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cab,
      DO(16) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cac,
      DO(15) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9d,
      DO(14) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9e,
      DO(13) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9f,
      DO(12) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca0,
      DO(11) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca1,
      DO(10) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca2,
      DO(9) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca3,
      DO(8) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca4,
      DO(7) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c95,
      DO(6) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c96,
      DO(5) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c97,
      DO(4) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c98,
      DO(3) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c99,
      DO(2) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9a,
      DO(1) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9b,
      DO(0) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9c,
      WRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007d7,
      WRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007d8,
      WRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007d9,
      WRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007da,
      WRADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      WRADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      WRADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      WRADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      WRADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      RDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007e4,
      RDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007e0,
      RDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007e5,
      RDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007e6,
      RDADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      RDADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      RDADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      RDADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      RDADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DI(31) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DI(30) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DI(29) => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5,
      DI(28) => blk00000001_blk000001a2_blk000001a3_sig000008a9,
      DI(27) => blk00000001_blk000001a2_blk000001a3_sig000008a8,
      DI(26) => blk00000001_blk000001a2_blk000001a3_sig000008a7,
      DI(25) => blk00000001_blk000001a2_blk000001a3_sig000008a6,
      DI(24) => blk00000001_blk000001a2_blk000001a3_sig000008a5,
      DI(23) => blk00000001_blk000001a2_blk000001a3_sig000008a3,
      DI(22) => blk00000001_blk000001a2_blk000001a3_sig000008a2,
      DI(21) => blk00000001_blk000001a2_blk000001a3_sig000008a1,
      DI(20) => blk00000001_blk000001a2_blk000001a3_sig000008a0,
      DI(19) => blk00000001_blk000001a2_blk000001a3_sig0000089f,
      DI(18) => blk00000001_blk000001a2_blk000001a3_sig0000089e,
      DI(17) => blk00000001_blk000001a2_blk000001a3_sig0000089d,
      DI(16) => blk00000001_blk000001a2_blk000001a3_sig0000089c,
      DI(15) => blk00000001_blk000001a2_blk000001a3_sig0000089a,
      DI(14) => blk00000001_blk000001a2_blk000001a3_sig00000899,
      DI(13) => blk00000001_blk000001a2_blk000001a3_sig00000898,
      DI(12) => blk00000001_blk000001a2_blk000001a3_sig00000897,
      DI(11) => blk00000001_blk000001a2_blk000001a3_sig00000896,
      DI(10) => blk00000001_blk000001a2_blk000001a3_sig00000895,
      DI(9) => blk00000001_blk000001a2_blk000001a3_sig00000894,
      DI(8) => blk00000001_blk000001a2_blk000001a3_sig00000893,
      DI(7) => blk00000001_blk000001a2_blk000001a3_sig00000891,
      DI(6) => blk00000001_blk000001a2_blk000001a3_sig00000890,
      DI(5) => blk00000001_blk000001a2_blk000001a3_sig0000088f,
      DI(4) => blk00000001_blk000001a2_blk000001a3_sig0000088e,
      DI(3) => blk00000001_blk000001a2_blk000001a3_sig0000088d,
      DI(2) => blk00000001_blk000001a2_blk000001a3_sig0000088c,
      DI(1) => blk00000001_blk000001a2_blk000001a3_sig0000088b,
      DI(0) => blk00000001_blk000001a2_blk000001a3_sig0000088a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d72 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cad,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000829
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d71 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cae,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000828
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d70 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caf,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000827
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000826
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000825
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000824
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000823
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000822
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d6a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000821
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d69 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000820
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d68 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca9,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d67 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001caa,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d66 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cab,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d65 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cac,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d64 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb3,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d63 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9d,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000081a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d62 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000819
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d61 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000818
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d60 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca0,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000817
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca1,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000816
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000815
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca3,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000814
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001ca4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000813
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cb2,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000812
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d5a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c95,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000811
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d59 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c96,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000810
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d58 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c97,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d57 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c98,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d56 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c99,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d55 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9a,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d54 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9b,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d53 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001c9c,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000080a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d51_blk00000d52 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000d51_sig00001cd5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000009a,
      RDCLK => aclk,
      WREN => blk00000001_sig0000009a,
      RDEN => blk00000001_sig0000009a,
      WRCLK => aclk,
      SSR => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DIP(3) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DIP(2) => blk00000001_blk000001a2_blk000001a3_sig000008c4,
      DIP(1) => blk00000001_blk000001a2_blk000001a3_sig000008bb,
      DIP(0) => blk00000001_blk000001a2_blk000001a3_sig000008b2,
      DOP(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d21,
      DOP(1) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d20,
      DOP(0) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1f,
      WE(3) => blk00000001_blk000001a2_blk000001a3_sig000007c9,
      WE(2) => blk00000001_blk000001a2_blk000001a3_sig000007c9,
      WE(1) => blk00000001_blk000001a2_blk000001a3_sig000007c9,
      WE(0) => blk00000001_blk000001a2_blk000001a3_sig000007c9,
      DO(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d96_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1a,
      DO(27) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1b,
      DO(26) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1c,
      DO(25) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1d,
      DO(24) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1e,
      DO(23) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d12,
      DO(22) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d13,
      DO(21) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d14,
      DO(20) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d15,
      DO(19) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d16,
      DO(18) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d17,
      DO(17) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d18,
      DO(16) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d19,
      DO(15) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0a,
      DO(14) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0b,
      DO(13) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0c,
      DO(12) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0d,
      DO(11) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0e,
      DO(10) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0f,
      DO(9) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d10,
      DO(8) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d11,
      DO(7) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d02,
      DO(6) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d03,
      DO(5) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d04,
      DO(4) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d05,
      DO(3) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d06,
      DO(2) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d07,
      DO(1) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d08,
      DO(0) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d09,
      WRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007d3,
      WRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007d4,
      WRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007d5,
      WRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007d6,
      WRADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      WRADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      WRADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      WRADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      WRADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      RDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007e2,
      RDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007dc,
      RDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007e3,
      RDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007de,
      RDADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      RDADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      RDADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      RDADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      RDADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DI(31) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DI(30) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DI(29) => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42,
      DI(28) => blk00000001_blk000001a2_blk000001a3_sig000008c9,
      DI(27) => blk00000001_blk000001a2_blk000001a3_sig000008c8,
      DI(26) => blk00000001_blk000001a2_blk000001a3_sig000008c7,
      DI(25) => blk00000001_blk000001a2_blk000001a3_sig000008c6,
      DI(24) => blk00000001_blk000001a2_blk000001a3_sig000008c5,
      DI(23) => blk00000001_blk000001a2_blk000001a3_sig000008c3,
      DI(22) => blk00000001_blk000001a2_blk000001a3_sig000008c2,
      DI(21) => blk00000001_blk000001a2_blk000001a3_sig000008c1,
      DI(20) => blk00000001_blk000001a2_blk000001a3_sig000008c0,
      DI(19) => blk00000001_blk000001a2_blk000001a3_sig000008bf,
      DI(18) => blk00000001_blk000001a2_blk000001a3_sig000008be,
      DI(17) => blk00000001_blk000001a2_blk000001a3_sig000008bd,
      DI(16) => blk00000001_blk000001a2_blk000001a3_sig000008bc,
      DI(15) => blk00000001_blk000001a2_blk000001a3_sig000008ba,
      DI(14) => blk00000001_blk000001a2_blk000001a3_sig000008b9,
      DI(13) => blk00000001_blk000001a2_blk000001a3_sig000008b8,
      DI(12) => blk00000001_blk000001a2_blk000001a3_sig000008b7,
      DI(11) => blk00000001_blk000001a2_blk000001a3_sig000008b6,
      DI(10) => blk00000001_blk000001a2_blk000001a3_sig000008b5,
      DI(9) => blk00000001_blk000001a2_blk000001a3_sig000008b4,
      DI(8) => blk00000001_blk000001a2_blk000001a3_sig000008b3,
      DI(7) => blk00000001_blk000001a2_blk000001a3_sig000008b1,
      DI(6) => blk00000001_blk000001a2_blk000001a3_sig000008b0,
      DI(5) => blk00000001_blk000001a2_blk000001a3_sig000008af,
      DI(4) => blk00000001_blk000001a2_blk000001a3_sig000008ae,
      DI(3) => blk00000001_blk000001a2_blk000001a3_sig000008ad,
      DI(2) => blk00000001_blk000001a2_blk000001a3_sig000008ac,
      DI(1) => blk00000001_blk000001a2_blk000001a3_sig000008ab,
      DI(0) => blk00000001_blk000001a2_blk000001a3_sig000008aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d95 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000849
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d94 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000848
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d93 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000847
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d92 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000846
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d91 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000845
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d90 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d21,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000844
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d12,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000843
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d13,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000842
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d14,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000841
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d15,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000840
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d16,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d8a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d17,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d89 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d18,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d88 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d19,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d87 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d20,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d86 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0a,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000083a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d85 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000839
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d84 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000838
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d83 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000837
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d82 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000836
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d81 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d0f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000835
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d80 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d10,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000834
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d11,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000833
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d1f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000832
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d02,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000831
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d03,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000830
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d04,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d7a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d05,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d79 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d06,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d78 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d07,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d77 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d08,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d76 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d09,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000082a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d74_blk00000d75 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000d74_sig00001d42
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9 : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000009a,
      RDCLK => aclk,
      WREN => blk00000001_sig0000009a,
      RDEN => blk00000001_sig0000009a,
      WRCLK => aclk,
      SSR => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DIP(3) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DIP(2) => blk00000001_blk000001a2_blk000001a3_sig000008e4,
      DIP(1) => blk00000001_blk000001a2_blk000001a3_sig000008db,
      DIP(0) => blk00000001_blk000001a2_blk000001a3_sig000008d2,
      DOP(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8e,
      DOP(1) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8d,
      DOP(0) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8c,
      WE(3) => blk00000001_blk000001a2_blk000001a3_sig000007c8,
      WE(2) => blk00000001_blk000001a2_blk000001a3_sig000007c8,
      WE(1) => blk00000001_blk000001a2_blk000001a3_sig000007c8,
      WE(0) => blk00000001_blk000001a2_blk000001a3_sig000007c8,
      DO(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db9_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d87,
      DO(27) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d88,
      DO(26) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d89,
      DO(25) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8a,
      DO(24) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8b,
      DO(23) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7f,
      DO(22) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d80,
      DO(21) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d81,
      DO(20) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d82,
      DO(19) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d83,
      DO(18) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d84,
      DO(17) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d85,
      DO(16) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d86,
      DO(15) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d77,
      DO(14) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d78,
      DO(13) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d79,
      DO(12) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7a,
      DO(11) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7b,
      DO(10) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7c,
      DO(9) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7d,
      DO(8) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7e,
      DO(7) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d6f,
      DO(6) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d70,
      DO(5) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d71,
      DO(4) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d72,
      DO(3) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d73,
      DO(2) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d74,
      DO(1) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d75,
      DO(0) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d76,
      WRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007cf,
      WRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007d0,
      WRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007d1,
      WRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007d2,
      WRADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      WRADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      WRADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      WRADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      WRADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      RDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007df,
      RDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007e0,
      RDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007e1,
      RDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007e6,
      RDADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      RDADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      RDADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      RDADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      RDADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DI(31) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DI(30) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DI(29) => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf,
      DI(28) => blk00000001_blk000001a2_blk000001a3_sig000008e9,
      DI(27) => blk00000001_blk000001a2_blk000001a3_sig000008e8,
      DI(26) => blk00000001_blk000001a2_blk000001a3_sig000008e7,
      DI(25) => blk00000001_blk000001a2_blk000001a3_sig000008e6,
      DI(24) => blk00000001_blk000001a2_blk000001a3_sig000008e5,
      DI(23) => blk00000001_blk000001a2_blk000001a3_sig000008e3,
      DI(22) => blk00000001_blk000001a2_blk000001a3_sig000008e2,
      DI(21) => blk00000001_blk000001a2_blk000001a3_sig000008e1,
      DI(20) => blk00000001_blk000001a2_blk000001a3_sig000008e0,
      DI(19) => blk00000001_blk000001a2_blk000001a3_sig000008df,
      DI(18) => blk00000001_blk000001a2_blk000001a3_sig000008de,
      DI(17) => blk00000001_blk000001a2_blk000001a3_sig000008dd,
      DI(16) => blk00000001_blk000001a2_blk000001a3_sig000008dc,
      DI(15) => blk00000001_blk000001a2_blk000001a3_sig000008da,
      DI(14) => blk00000001_blk000001a2_blk000001a3_sig000008d9,
      DI(13) => blk00000001_blk000001a2_blk000001a3_sig000008d8,
      DI(12) => blk00000001_blk000001a2_blk000001a3_sig000008d7,
      DI(11) => blk00000001_blk000001a2_blk000001a3_sig000008d6,
      DI(10) => blk00000001_blk000001a2_blk000001a3_sig000008d5,
      DI(9) => blk00000001_blk000001a2_blk000001a3_sig000008d4,
      DI(8) => blk00000001_blk000001a2_blk000001a3_sig000008d3,
      DI(7) => blk00000001_blk000001a2_blk000001a3_sig000008d1,
      DI(6) => blk00000001_blk000001a2_blk000001a3_sig000008d0,
      DI(5) => blk00000001_blk000001a2_blk000001a3_sig000008cf,
      DI(4) => blk00000001_blk000001a2_blk000001a3_sig000008ce,
      DI(3) => blk00000001_blk000001a2_blk000001a3_sig000008cd,
      DI(2) => blk00000001_blk000001a2_blk000001a3_sig000008cc,
      DI(1) => blk00000001_blk000001a2_blk000001a3_sig000008cb,
      DI(0) => blk00000001_blk000001a2_blk000001a3_sig000008ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d87,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000869
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d88,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000868
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d89,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000867
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000866
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000865
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000864
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000863
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d80,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000862
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000db0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d81,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000861
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000daf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d82,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000860
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000dae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d83,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000dad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d84,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000dac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d85,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000dab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d86,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000daa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8d,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d77,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000085a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d78,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000859
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d79,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000858
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000857
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000856
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000855
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7d,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000854
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d7e,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000853
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d8c,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000852
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000da0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d6f,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000851
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d70,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000850
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d71,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d72,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d73,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d74,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d9a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d75,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d99 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001d76,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000084a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000d97_blk00000d98 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000d97_sig00001daf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc : RAMB18SDP
    generic map(
      DO_REG => 1,
      INIT => X"000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "GENERATE_X_ONLY",
      SIM_MODE => "SAFE",
      SRVAL => X"000000000"
    )
    port map (
      REGCE => blk00000001_sig0000009a,
      RDCLK => aclk,
      WREN => blk00000001_sig0000009a,
      RDEN => blk00000001_sig0000009a,
      WRCLK => aclk,
      SSR => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DIP(3) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DIP(2) => blk00000001_blk000001a2_blk000001a3_sig00000904,
      DIP(1) => blk00000001_blk000001a2_blk000001a3_sig000008fb,
      DIP(0) => blk00000001_blk000001a2_blk000001a3_sig000008f2,
      DOP(3) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DOP_3_UNCONNECTED,
      DOP(2) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfb,
      DOP(1) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfa,
      DOP(0) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df9,
      WE(3) => blk00000001_blk000001a2_blk000001a3_sig000007c7,
      WE(2) => blk00000001_blk000001a2_blk000001a3_sig000007c7,
      WE(1) => blk00000001_blk000001a2_blk000001a3_sig000007c7,
      WE(0) => blk00000001_blk000001a2_blk000001a3_sig000007c7,
      DO(31) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_31_UNCONNECTED,
      DO(30) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_30_UNCONNECTED,
      DO(29) => NLW_blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddc_DO_29_UNCONNECTED,
      DO(28) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df4,
      DO(27) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df5,
      DO(26) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df6,
      DO(25) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df7,
      DO(24) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df8,
      DO(23) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dec,
      DO(22) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ded,
      DO(21) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dee,
      DO(20) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001def,
      DO(19) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df0,
      DO(18) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df1,
      DO(17) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df2,
      DO(16) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df3,
      DO(15) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de4,
      DO(14) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de5,
      DO(13) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de6,
      DO(12) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de7,
      DO(11) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de8,
      DO(10) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de9,
      DO(9) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dea,
      DO(8) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001deb,
      DO(7) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddc,
      DO(6) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddd,
      DO(5) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dde,
      DO(4) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddf,
      DO(3) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de0,
      DO(2) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de1,
      DO(1) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de2,
      DO(0) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de3,
      WRADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007cb,
      WRADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007cc,
      WRADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007cd,
      WRADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007ce,
      WRADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      WRADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      WRADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      WRADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      WRADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      RDADDR(8) => blk00000001_blk000001a2_blk000001a3_sig000007db,
      RDADDR(7) => blk00000001_blk000001a2_blk000001a3_sig000007dc,
      RDADDR(6) => blk00000001_blk000001a2_blk000001a3_sig000007dd,
      RDADDR(5) => blk00000001_blk000001a2_blk000001a3_sig000007de,
      RDADDR(4) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      RDADDR(3) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      RDADDR(2) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      RDADDR(1) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      RDADDR(0) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DI(31) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DI(30) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DI(29) => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c,
      DI(28) => blk00000001_blk000001a2_blk000001a3_sig00000909,
      DI(27) => blk00000001_blk000001a2_blk000001a3_sig00000908,
      DI(26) => blk00000001_blk000001a2_blk000001a3_sig00000907,
      DI(25) => blk00000001_blk000001a2_blk000001a3_sig00000906,
      DI(24) => blk00000001_blk000001a2_blk000001a3_sig00000905,
      DI(23) => blk00000001_blk000001a2_blk000001a3_sig00000903,
      DI(22) => blk00000001_blk000001a2_blk000001a3_sig00000902,
      DI(21) => blk00000001_blk000001a2_blk000001a3_sig00000901,
      DI(20) => blk00000001_blk000001a2_blk000001a3_sig00000900,
      DI(19) => blk00000001_blk000001a2_blk000001a3_sig000008ff,
      DI(18) => blk00000001_blk000001a2_blk000001a3_sig000008fe,
      DI(17) => blk00000001_blk000001a2_blk000001a3_sig000008fd,
      DI(16) => blk00000001_blk000001a2_blk000001a3_sig000008fc,
      DI(15) => blk00000001_blk000001a2_blk000001a3_sig000008fa,
      DI(14) => blk00000001_blk000001a2_blk000001a3_sig000008f9,
      DI(13) => blk00000001_blk000001a2_blk000001a3_sig000008f8,
      DI(12) => blk00000001_blk000001a2_blk000001a3_sig000008f7,
      DI(11) => blk00000001_blk000001a2_blk000001a3_sig000008f6,
      DI(10) => blk00000001_blk000001a2_blk000001a3_sig000008f5,
      DI(9) => blk00000001_blk000001a2_blk000001a3_sig000008f4,
      DI(8) => blk00000001_blk000001a2_blk000001a3_sig000008f3,
      DI(7) => blk00000001_blk000001a2_blk000001a3_sig000008f1,
      DI(6) => blk00000001_blk000001a2_blk000001a3_sig000008f0,
      DI(5) => blk00000001_blk000001a2_blk000001a3_sig000008ef,
      DI(4) => blk00000001_blk000001a2_blk000001a3_sig000008ee,
      DI(3) => blk00000001_blk000001a2_blk000001a3_sig000008ed,
      DI(2) => blk00000001_blk000001a2_blk000001a3_sig000008ec,
      DI(1) => blk00000001_blk000001a2_blk000001a3_sig000008eb,
      DI(0) => blk00000001_blk000001a2_blk000001a3_sig000008ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000ddb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df4,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000889
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dda : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000888
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000887
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000886
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000885
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000884
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dec,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000883
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ded,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000882
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dee,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000881
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001def,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000880
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df0,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dd0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dcf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df2,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df3,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dcd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dfa,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dcc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de4,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000087a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dcb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de5,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000879
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de6,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000878
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de7,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000877
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de8,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000876
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000875
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dea,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000874
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001deb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000873
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001df9,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000872
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddc,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000871
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddd,
      Q => blk00000001_blk000001a2_blk000001a3_sig00000870
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001dde,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dc0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001ddf,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dbf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de0,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dbe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de1,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dbd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de2,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dbc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001de3,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000086a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000dba_blk00000dbb : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000dba_sig00001e1c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000de2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e28,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000de1 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e27,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e26,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e26,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e26,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000007fe,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e28,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000de1_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000de0 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e27
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_blk00000ddf : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ddd_blk00000dde_sig00001e26
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e34,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ea
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de7 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e33,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e32,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e32,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e32,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011eb,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e34,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de7_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de6 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e33
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_blk00000de5 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000de3_blk00000de4_sig00001e32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000dee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e40,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ec
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000ded : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3f,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3e,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3e,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3e,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e40,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000ded_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000dec : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_blk00000deb : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000de9_blk00000dea_sig00001e3e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4c,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df3 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4b,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4a,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4a,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4a,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig000000c7,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4c,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df3_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df2 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_blk00000df1 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000def_blk00000df0_sig00001e4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000dfa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e58,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007f5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000df9 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e57,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e56,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e56,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e56,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_sig000000c7,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e58,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000df9_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000df8 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_blk00000df7 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000df5_blk00000df6_sig00001e56
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e59 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001273,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e58 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001274,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e70
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e57 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001275,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e56 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001276,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e55 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001277,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e54 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e65,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e53 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6c,
      O => blk00000001_blk000001a2_blk000001a3_sig0000126c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e52 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e67,
      LI => blk00000001_blk000001a2_blk000001a3_sig00001278,
      O => blk00000001_blk000001a2_blk000001a3_sig00001271
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e51 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6b,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e70,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e50 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e70,
      O => blk00000001_blk000001a2_blk000001a3_sig0000126d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4f : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6a,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e69
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4e : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6f,
      O => blk00000001_blk000001a2_blk000001a3_sig0000126e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4d : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e69,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e68
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4c : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e69,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6e,
      O => blk00000001_blk000001a2_blk000001a3_sig0000126f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e68,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e67
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e4a : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e68,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e6d,
      O => blk00000001_blk000001a2_blk000001a3_sig00001270
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e49 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e66
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e47_blk00000e48 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000e47_sig00001e65
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e8d : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig0000128e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e87
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e8c : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig0000128f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e8b : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001290,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e8a : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001291,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e89 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001292,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e89
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e88 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001293,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e88
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e87 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e7f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e87,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e86
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e86 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e87,
      O => blk00000001_blk000001a2_blk000001a3_sig00001281
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e85 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e81,
      LI => blk00000001_blk000001a2_blk000001a3_sig00001294,
      O => blk00000001_blk000001a2_blk000001a3_sig00001287
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e84 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e86,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e85
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e83 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e86,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8c,
      O => blk00000001_blk000001a2_blk000001a3_sig00001282
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e82 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e85,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e84
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e81 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e85,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8b,
      O => blk00000001_blk000001a2_blk000001a3_sig00001283
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e80 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e84,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e83
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e84,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e8a,
      O => blk00000001_blk000001a2_blk000001a3_sig00001284
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e83,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e89,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e82
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e83,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e89,
      O => blk00000001_blk000001a2_blk000001a3_sig00001285
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e82,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e88,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e81
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e82,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e88,
      O => blk00000001_blk000001a2_blk000001a3_sig00001286
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e7a : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e80
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e78_blk00000e79 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000e78_sig00001e7f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000ea4 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig000012ac,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000ea3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012ad,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000ea2 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012ae,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000ea1 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e95,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9a,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e99
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000ea0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9a,
      O => blk00000001_blk000001a2_blk000001a3_sig000012a7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9f : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e97,
      LI => blk00000001_blk000001a2_blk000001a3_sig000012af,
      O => blk00000001_blk000001a2_blk000001a3_sig000012aa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9e : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e99,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e98
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9d : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e99,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9c,
      O => blk00000001_blk000001a2_blk000001a3_sig000012a8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9c : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e98,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96,
      S => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9b,
      O => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e97
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9b : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e98,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e9b,
      O => blk00000001_blk000001a2_blk000001a3_sig000012a9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e9a : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e96
    );
  blk00000001_blk000001a2_blk000001a3_blk00000e98_blk00000e99 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000e98_sig00001e95
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ec0 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig000012ba,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ead
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ebf : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012bb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eb0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ebe : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012bc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaf
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ebd : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012bd,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eae
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ebc : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea7,
      S => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ead,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eac
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000ebb : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ead,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eba : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea9,
      LI => blk00000001_blk000001a2_blk000001a3_sig000012be,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eac,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8,
      S => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eb0,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eab
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb8 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eac,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eb0,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eab,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8,
      S => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaf,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eab,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaf,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb5 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaa,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8,
      S => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eae,
      O => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eaa,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001eae,
      O => blk00000001_blk000001a2_blk000001a3_sig000012b7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb3 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eb1_blk00000eb2 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000eb1_sig00001ea7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001ebb,
      Q => blk00000001_blk000001a2_blk000001a3_sig0000124c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eba,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eb9,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eba,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eb9,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00001247,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001ebb,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec5_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec4 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eba
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_blk00000ec3 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ec1_blk00000ec2_sig00001eb9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ed4 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig000012cb,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ed3 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig000012cc,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ed2 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec3,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec2,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec6,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ed1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec3,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec6,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ed0 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec4,
      LI => blk00000001_blk000001a2_blk000001a3_sig000012cd,
      O => blk00000001_blk000001a2_blk000001a3_sig000012ca
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ecf : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec5,
      DI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec3,
      S => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec7,
      O => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ece : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec5,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec7,
      O => blk00000001_blk000001a2_blk000001a3_sig000012c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ecd : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec3
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ecb_blk00000ecc : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ecb_sig00001ec2
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000eda : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001edb,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001249
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000ed9 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig0000124a,
      CE => blk00000001_sig0000009a,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001edb,
      Q31 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000ed9_Q31_UNCONNECTED,
      A(4) => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001eda,
      A(3) => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9,
      A(2) => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9,
      A(1) => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9,
      A(0) => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000ed8 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001eda
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_blk00000ed7 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ed5_blk00000ed6_sig00001ed9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000ee0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee6,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011f6
    );
  blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000edf : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee4,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee4,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee5,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee4,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee6,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000edf_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000ede : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee5
    );
  blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_blk00000edd : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000edb_blk00000edc_sig00001ee4
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef1,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007f7
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee5 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef0,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef0,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001eef,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef0,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000801,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef1,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee5_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee4 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001ef0
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_blk00000ee3 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ee1_blk00000ee2_sig00001eef
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000eec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efc,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007f8
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000eeb : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efa,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efb,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efb,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efb,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig00000801,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efc,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000eeb_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000eea : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_blk00000ee9 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ee7_blk00000ee8_sig00001efa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000ef2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f10,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007fa
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000ef1 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      CE => blk00000001_sig0000009a,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f10,
      Q31 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000ef1_Q31_UNCONNECTED,
      A(4) => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0f,
      A(3) => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e,
      A(2) => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e,
      A(1) => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e,
      A(0) => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000ef0 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_blk00000eef : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000eed_blk00000eee_sig00001f0e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f24,
      Q => blk00000001_blk000001a2_blk000001a3_sig000007fb
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef7 : SRLC32E
    generic map(
      INIT => X"00000000"
    )
    port map (
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fb,
      CE => blk00000001_sig0000009a,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f24,
      Q31 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef7_Q31_UNCONNECTED,
      A(4) => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f23,
      A(3) => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22,
      A(2) => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22,
      A(1) => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22,
      A(0) => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef6 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f23
    );
  blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_blk00000ef5 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000ef3_blk00000ef4_sig00001f22
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f19 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f32,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f2f,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f19_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f18 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      Q => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f18_Q_UNCONNECTED,
      Q15 => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f32
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f17 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f31
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f16 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f30
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_blk00000f15 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f13_blk00000f14_sig00001f2f,
      R => blk00000001_blk000001a2_blk000001a3_sig000011f7,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ee
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3d,
      Q => blk00000001_blk000001a2_blk000001a3_sig000011ed
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1e : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3b,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3c,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3c,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3b,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011f9,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3d,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1e_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1d : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_blk00000f1c : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000f1a_blk00000f1b_sig00001f3b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f25 : SRLC16E
    generic map(
      INIT => X"0000"
    )
    port map (
      A0 => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f49,
      A1 => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f4a,
      A2 => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f4a,
      A3 => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f49,
      CE => blk00000001_sig0000009a,
      CLK => aclk,
      D => blk00000001_blk000001a2_blk000001a3_sig000011fa,
      Q => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f48,
      Q15 => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f25_Q15_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f24 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f4a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f23 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f49
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_blk00000f22 : FDRE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f20_blk00000f21_sig00001f48,
      R => blk00000001_blk000001a2_blk000001a3_sig000007f9,
      Q => blk00000001_sig000000c9
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f64 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001311,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5f
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f63 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig00001310,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f62 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig0000130f,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f61 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig0000130e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f60 : INV
    port map (
      I => blk00000001_blk000001a2_blk000001a3_sig0000130e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f60
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f58,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001301
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5b,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001302
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5a,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001303
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => aclk,
      CE => blk00000001_sig0000009a,
      D => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f59,
      Q => blk00000001_blk000001a2_blk000001a3_sig00001304
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5b : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f57,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f60,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f64
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f5a : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f64,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000130e,
      S => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f63
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f59 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f63,
      DI => blk00000001_blk000001a2_blk000001a3_sig0000130f,
      S => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f62
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f58 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f62,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001310,
      S => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f61
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f57 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f64,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f56 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f63,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f55 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f62,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5c,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f59
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f54 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f61,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f5f,
      O => NLW_blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f54_O_UNCONNECTED
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f53 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f57,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f60,
      O => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f58
    );
  blk00000001_blk000001a2_blk000001a3_blk00000f51_blk00000f52 : VCC
    port map (
      P => blk00000001_blk000001a2_blk000001a3_blk00000f51_sig00001f57
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00001000 : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001354,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7e
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000fff : LUT1
    generic map(
      INIT => X"2"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001351,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7d
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ffe : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001351,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001352,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f75
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ffd : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001352,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001353,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f76
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ffc : LUT2
    generic map(
      INIT => X"6"
    )
    port map (
      I0 => blk00000001_blk000001a2_blk000001a3_sig00001353,
      I1 => blk00000001_blk000001a2_blk000001a3_sig00001354,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f77
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ffb : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f74,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001354,
      S => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7e,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7c
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ffa : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7c,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001353,
      S => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f77,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7b
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff9 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7b,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001352,
      S => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f76,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff8 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7a,
      DI => blk00000001_blk000001a2_blk000001a3_sig00001351,
      S => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f75,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f79
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff7 : MUXCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f79,
      DI => blk00000001_blk000001a2_sig00000592,
      S => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7d,
      O => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f78
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff6 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7c,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f77,
      O => blk00000001_blk000001a2_blk000001a3_sig00001356
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff5 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7b,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f76,
      O => blk00000001_blk000001a2_blk000001a3_sig00001357
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff4 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7a,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f75,
      O => blk00000001_blk000001a2_blk000001a3_sig00001358
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff3 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f79,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7d,
      O => blk00000001_blk000001a2_blk000001a3_sig00001359
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff2 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f78,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f74,
      O => blk00000001_blk000001a2_blk000001a3_sig0000135a
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff1 : XORCY
    port map (
      CI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f74,
      LI => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f7e,
      O => blk00000001_blk000001a2_blk000001a3_sig00001355
    );
  blk00000001_blk000001a2_blk000001a3_blk00000fef_blk00000ff0 : GND
    port map (
      G => blk00000001_blk000001a2_blk000001a3_blk00000fef_sig00001f74
    );

end STRUCTURE;

-- synthesis translate_on

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlFloat : integer := 3;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function shift_division_result(quotient, fraction: std_logic_vector;
                                   fraction_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant q_width : integer := quotient'length;
        constant f_width : integer := fraction'length;
        constant vec_MSB : integer := q_width+f_width-1;
        constant result_MSB : integer := q_width+fraction_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := ( quotient & fraction );
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function shift_op (inp: std_logic_vector;
                       result_width, shift_value, shift_dir: INTEGER)
        return std_logic_vector
    is
        constant inp_width : integer := inp'length;
        constant vec_MSB : integer := inp_width-1;
        constant result_MSB : integer := result_width-1;
        constant result_LSB : integer := vec_MSB-result_MSB;
        variable vec : std_logic_vector(vec_MSB downto 0);
        variable result : std_logic_vector(result_MSB downto 0);
    begin
        vec := inp;
        if shift_dir = 1 then
            for i in vec_MSB downto 0 loop
                if (i < shift_value) then
                     vec(i) := '0';
                else
                    vec(i) := vec(i-shift_value);
                end if;
            end loop;
        else
            for i in 0 to vec_MSB loop
                if (i > vec_MSB-shift_value) then
                    vec(i) := vec(vec_MSB);
                else
                    vec(i) := vec(i+shift_value);
                end if;
            end loop;
        end if;
        result := vec(vec_MSB downto result_LSB);
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if clr = '1' then
            reg_bank_in <= (others => (others => '0'));
          elsif ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlclockenablegenerator is
  generic (
    period: integer := 2;
    log_2_period: integer := 0;
    pipeline_regs: integer := 5
  );
  port (
    clk: in std_logic;
    clr: in std_logic;
    ce: out std_logic
  );
end xlclockenablegenerator;
architecture behavior of xlclockenablegenerator is
  component synth_reg_w_init
    generic (
      width: integer;
      init_index: integer;
      init_value: bit_vector;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function size_of_uint(inp: integer; power_of_2: boolean)
    return integer
  is
    constant inp_vec: std_logic_vector(31 downto 0) :=
      integer_to_std_logic_vector(inp,32, xlUnsigned);
    variable result: integer;
  begin
    result := 32;
    for i in 0 to 31 loop
      if inp_vec(i) = '1' then
        result := i;
      end if;
    end loop;
    if power_of_2 then
      return result;
    else
      return result+1;
    end if;
  end;
  function is_power_of_2(inp: std_logic_vector)
    return boolean
  is
    constant width: integer := inp'length;
    variable vec: std_logic_vector(width - 1 downto 0);
    variable single_bit_set: boolean;
    variable more_than_one_bit_set: boolean;
    variable result: boolean;
  begin
    vec := inp;
    single_bit_set := false;
    more_than_one_bit_set := false;
    -- synopsys translate_off
    if (is_XorU(vec)) then
      return false;
    end if;
     -- synopsys translate_on
    if width > 0 then
      for i in 0 to width - 1 loop
        if vec(i) = '1' then
          if single_bit_set then
            more_than_one_bit_set := true;
          end if;
          single_bit_set := true;
        end if;
      end loop;
    end if;
    if (single_bit_set and not(more_than_one_bit_set)) then
      result := true;
    else
      result := false;
    end if;
    return result;
  end;
  function ce_reg_init_val(index, period : integer)
    return integer
  is
     variable result: integer;
   begin
      result := 0;
      if ((index mod period) = 0) then
          result := 1;
      end if;
      return result;
  end;
  function remaining_pipe_regs(num_pipeline_regs, period : integer)
    return integer
  is
     variable factor, result: integer;
  begin
      factor := (num_pipeline_regs / period);
      result := num_pipeline_regs - (period * factor) + 1;
      return result;
  end;

  function sg_min(L, R: INTEGER) return INTEGER is
  begin
      if L < R then
            return L;
      else
            return R;
      end if;
  end;
  constant max_pipeline_regs : integer := 8;
  constant pipe_regs : integer := 5;
  constant num_pipeline_regs : integer := sg_min(pipeline_regs, max_pipeline_regs);
  constant rem_pipeline_regs : integer := remaining_pipe_regs(num_pipeline_regs,period);
  constant period_floor: integer := max(2, period);
  constant power_of_2_counter: boolean :=
    is_power_of_2(integer_to_std_logic_vector(period_floor,32, xlUnsigned));
  constant cnt_width: integer :=
    size_of_uint(period_floor, power_of_2_counter);
  constant clk_for_ce_pulse_minus1: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector((period_floor - 2),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus2: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - 3),cnt_width, xlUnsigned);
  constant clk_for_ce_pulse_minus_regs: std_logic_vector(cnt_width - 1 downto 0) :=
    integer_to_std_logic_vector(max(0,period - rem_pipeline_regs),cnt_width, xlUnsigned);
  signal clk_num: unsigned(cnt_width - 1 downto 0) := (others => '0');
  signal ce_vec : std_logic_vector(num_pipeline_regs downto 0);
  signal internal_ce: std_logic_vector(0 downto 0);
  signal cnt_clr, cnt_clr_dly: std_logic_vector (0 downto 0);
begin
  cntr_gen: process(clk)
  begin
    if clk'event and clk = '1'  then
        if ((cnt_clr_dly(0) = '1') or (clr = '1')) then
          clk_num <= (others => '0');
        else
          clk_num <= clk_num + 1;
        end if;
    end if;
  end process;
  clr_gen: process(clk_num, clr)
  begin
    if power_of_2_counter then
      cnt_clr(0) <= clr;
    else
      if (unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus1
          or clr = '1') then
        cnt_clr(0) <= '1';
      else
        cnt_clr(0) <= '0';
      end if;
    end if;
  end process;
  clr_reg: synth_reg_w_init
    generic map (
      width => 1,
      init_index => 0,
      init_value => b"0000",
      latency => 1
    )
    port map (
      i => cnt_clr,
      ce => '1',
      clr => clr,
      clk => clk,
      o => cnt_clr_dly
    );
  pipelined_ce : if period > 1 generate
      ce_gen: process(clk_num)
      begin
          if unsigned_to_std_logic_vector(clk_num) = clk_for_ce_pulse_minus_regs then
              ce_vec(num_pipeline_regs) <= '1';
          else
              ce_vec(num_pipeline_regs) <= '0';
          end if;
      end process;
      ce_pipeline: for index in num_pipeline_regs downto 1 generate
          ce_reg : synth_reg_w_init
              generic map (
                  width => 1,
                  init_index => ce_reg_init_val(index, period),
                  init_value => b"0000",
                  latency => 1
                  )
              port map (
                  i => ce_vec(index downto index),
                  ce => '1',
                  clr => clr,
                  clk => clk,
                  o => ce_vec(index-1 downto index-1)
                  );
      end generate;
      internal_ce <= ce_vec(0 downto 0);
  end generate;
  generate_clock_enable: if period > 1 generate
    ce <= internal_ce(0);
  end generate;
  generate_clock_enable_constant: if period = 1 generate
    ce <= '1';
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity accum_a764547d38 is
  port (
    b : in std_logic_vector((5 - 1) downto 0);
    rst : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((15 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end accum_a764547d38;


architecture behavior of accum_a764547d38 is
  signal b_17_24: unsigned((5 - 1) downto 0);
  signal rst_17_27: boolean;
  signal en_17_32: boolean;
  signal accum_reg_41_23: unsigned((15 - 1) downto 0) := "000000000000000";
  signal accum_reg_41_23_rst: std_logic;
  signal accum_reg_41_23_en: std_logic;
  signal cast_51_42: unsigned((15 - 1) downto 0);
  signal accum_reg_join_47_1: unsigned((16 - 1) downto 0);
  signal accum_reg_join_47_1_en: std_logic;
  signal accum_reg_join_47_1_rst: std_logic;
begin
  b_17_24 <= std_logic_vector_to_unsigned(b);
  rst_17_27 <= ((rst) = "1");
  en_17_32 <= ((en) = "1");
  proc_accum_reg_41_23: process (clk)
  is
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (accum_reg_41_23_rst = '1')) then
        accum_reg_41_23 <= "000000000000000";
      elsif ((ce = '1') and (accum_reg_41_23_en = '1')) then 
        accum_reg_41_23 <= accum_reg_41_23 + cast_51_42;
      end if;
    end if;
  end process proc_accum_reg_41_23;
  cast_51_42 <= u2u_cast(b_17_24, 0, 15, 0);
  proc_if_47_1: process (accum_reg_41_23, cast_51_42, en_17_32, rst_17_27)
  is
  begin
    if rst_17_27 then
      accum_reg_join_47_1_rst <= '1';
    elsif en_17_32 then
      accum_reg_join_47_1_rst <= '0';
    else 
      accum_reg_join_47_1_rst <= '0';
    end if;
    if en_17_32 then
      accum_reg_join_47_1_en <= '1';
    else 
      accum_reg_join_47_1_en <= '0';
    end if;
  end process proc_if_47_1;
  accum_reg_41_23_rst <= accum_reg_join_47_1_rst;
  accum_reg_41_23_en <= accum_reg_join_47_1_en;
  q <= unsigned_to_std_logic_vector(accum_reg_41_23);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xladdsub_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub_wlan_phy_tx_pmd;
architecture behavior of xladdsub_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_913f4bce6842c815
    port (
          a: in std_logic_vector(13 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(13 - 1 downto 0)
    );
  end component;
  component addsb_11_0_73986f767e994888
    port (
          a: in std_logic_vector(10 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(10 - 1 downto 0)
    );
  end component;
  component addsb_11_0_8dc9188fad4d9a9c
    port (
          a: in std_logic_vector(9 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(9 - 1 downto 0)
    );
  end component;
  component addsb_11_0_a52ead9b8a3c1e76
    port (
          a: in std_logic_vector(9 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(9 - 1 downto 0)
    );
  end component;
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_913f4bce6842c815")) generate
    core_instance0: addsb_11_0_913f4bce6842c815
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp2: if ((core_name0 = "addsb_11_0_73986f767e994888")) generate
    core_instance2: addsb_11_0_73986f767e994888
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp3: if ((core_name0 = "addsb_11_0_8dc9188fad4d9a9c")) generate
    core_instance3: addsb_11_0_8dc9188fad4d9a9c
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  comp4: if ((core_name0 = "addsb_11_0_a52ead9b8a3c1e76")) generate
    core_instance4: addsb_11_0_a52ead9b8a3c1e76
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlpassthrough is
    generic (
        din_width    : integer := 16;
        dout_width   : integer := 16
        );
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlpassthrough;
architecture passthrough_arch of xlpassthrough is
begin
  dout <= din;
end passthrough_arch;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlslice is
    generic (
        new_msb      : integer := 9;
        new_lsb      : integer := 1;
        x_width      : integer := 16;
        y_width      : integer := 8);
    port (
        x : in std_logic_vector (x_width-1 downto 0);
        y : out std_logic_vector (y_width-1 downto 0));
end xlslice;
architecture behavior of xlslice is
begin
    y <= x(new_msb downto new_lsb);
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_32afb77cd2 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_32afb77cd2;


architecture behavior of concat_32afb77cd2 is
  signal in0_1_23: boolean;
  signal in1_1_27: boolean;
  signal y_2_1_concat: unsigned((2 - 1) downto 0);
begin
  in0_1_23 <= ((in0) = "1");
  in1_1_27 <= ((in1) = "1");
  y_2_1_concat <= std_logic_vector_to_unsigned(boolean_to_vector(in0_1_23) & boolean_to_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a7e2bb9e12 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a7e2bb9e12;


architecture behavior of constant_a7e2bb9e12 is
begin
  op <= "01";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_a629aefb53 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a629aefb53;


architecture behavior of constant_a629aefb53 is
begin
  op <= "1001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_f5633478bf is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_f5633478bf;


architecture behavior of constant_f5633478bf is
begin
  op <= "10001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_07db25d611 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_07db25d611;


architecture behavior of constant_07db25d611 is
begin
  op <= "10111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_ef95fb0eb4 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_ef95fb0eb4;


architecture behavior of constant_ef95fb0eb4 is
begin
  op <= "101111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_145086465d is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_145086465d;


architecture behavior of constant_145086465d is
begin
  op <= "1000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_bc74ae1a6c is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_bc74ae1a6c;


architecture behavior of constant_bc74ae1a6c is
begin
  op <= "11000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_469094441c is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_469094441c;


architecture behavior of constant_469094441c is
begin
  op <= "100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4e64dfaf34 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4e64dfaf34;


architecture behavior of constant_4e64dfaf34 is
begin
  op <= "101";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer :=  0;
           reset        : integer :=  0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        rst     : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if ((reg_retiming = 0) and (reset = 0)) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if ((reg_retiming = 1) or (reset = 1)) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => rst,
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e5b38cca3b is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e5b38cca3b;


architecture behavior of inverter_e5b38cca3b is
  signal ip_1_26: boolean;
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of boolean;
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => false);
  signal op_mem_22_20_front_din: boolean;
  signal op_mem_22_20_back: boolean;
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: boolean;
begin
  ip_1_26 <= ((ip) = "1");
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= ((not boolean_to_vector(ip_1_26)) = "1");
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= boolean_to_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_80f90b97d0 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_80f90b97d0;


architecture behavior of logical_80f90b97d0 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_954ee29728 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_954ee29728;


architecture behavior of logical_954ee29728 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  fully_2_1_bit <= d0_1_24 and d1_1_27 and d2_1_30;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4a20039e59 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((4 - 1) downto 0);
    d2 : in std_logic_vector((5 - 1) downto 0);
    y : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4a20039e59;


architecture behavior of mux_4a20039e59 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((4 - 1) downto 0);
  signal d2_1_30: std_logic_vector((5 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((5 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 5, 0, xlUnsigned);
      when "01" =>
        unregy_join_6_1 <= cast(d1_1_27, 0, 5, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_ec1b27521c is
  port (
    a : in std_logic_vector((15 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_ec1b27521c;


architecture behavior of relational_ec1b27521c is
  signal a_1_31: unsigned((15 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal cast_12_17: unsigned((15 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 15, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_37ecee0ab7 is
  port (
    a : in std_logic_vector((15 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_37ecee0ab7;


architecture behavior of relational_37ecee0ab7 is
  signal a_1_31: unsigned((15 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal cast_12_17: unsigned((15 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 15, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_eed86727d9 is
  port (
    a : in std_logic_vector((15 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_eed86727d9;


architecture behavior of relational_eed86727d9 is
  signal a_1_31: unsigned((15 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal cast_16_16: unsigned((15 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_16_16 <= u2u_cast(b_1_34, 0, 15, 0);
  result_16_3_rel <= a_1_31 < cast_16_16;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_70fbe7d900 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_70fbe7d900;


architecture behavior of relational_70fbe7d900 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_b307c14bb5 is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_b307c14bb5;


architecture behavior of relational_b307c14bb5 is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_22_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_22_3_rel <= a_1_31 >= b_1_34;
  op <= boolean_to_vector(result_22_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_07bde14ec5 is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_07bde14ec5;


architecture behavior of relational_07bde14ec5 is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;
entity xlcounter_limit_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned;
    cnt_63_48: integer:= 0;
    cnt_47_32: integer:= 0;
    cnt_31_16: integer:= 0;
    cnt_15_0: integer:= 0;
    count_limited: integer := 0
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_limit_wlan_phy_tx_pmd ;
architecture behavior of xlcounter_limit_wlan_phy_tx_pmd is
  signal high_cnt_to: std_logic_vector(31 downto 0);
  signal low_cnt_to: std_logic_vector(31 downto 0);
  signal cnt_to: std_logic_vector(63 downto 0);
  signal core_sinit, op_thresh0, core_ce: std_logic;
  signal rst_overrides_en: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
  -- synopsys translate_off
  signal real_op : real;
   -- synopsys translate_on
  function equals(op, cnt_to : std_logic_vector; width, arith : integer)
    return std_logic
  is
    variable signed_op, signed_cnt_to : signed (width - 1 downto 0);
    variable unsigned_op, unsigned_cnt_to : unsigned (width - 1 downto 0);
    variable result : std_logic;
  begin
    -- synopsys translate_off
    if ((is_XorU(op)) or (is_XorU(cnt_to)) ) then
      result := '0';
      return result;
    end if;
    -- synopsys translate_on
    if (op = cnt_to) then
      result := '1';
    else
      result := '0';
    end if;
    return result;
  end;
  component cntr_11_0_bcc28bfecf25caff
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_bcc28bfecf25caff:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_bcc28bfecf25caff:
    component is "true";
  attribute box_type of cntr_11_0_bcc28bfecf25caff:
    component  is "black_box";
  component cntr_11_0_86806e294f737f4c
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_86806e294f737f4c:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_86806e294f737f4c:
    component is "true";
  attribute box_type of cntr_11_0_86806e294f737f4c:
    component  is "black_box";
  component cntr_11_0_36e2bb554c95560d
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_36e2bb554c95560d:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_36e2bb554c95560d:
    component is "true";
  attribute box_type of cntr_11_0_36e2bb554c95560d:
    component  is "black_box";
  component cntr_11_0_f068fb73312ae1e5
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_f068fb73312ae1e5:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_f068fb73312ae1e5:
    component is "true";
  attribute box_type of cntr_11_0_f068fb73312ae1e5:
    component  is "black_box";
  component cntr_11_0_d24951bef2f0cdc9
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d24951bef2f0cdc9:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d24951bef2f0cdc9:
    component is "true";
  attribute box_type of cntr_11_0_d24951bef2f0cdc9:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec : std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec : std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr : string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
begin
  -- synopsys translate_off
  -- synopsys translate_on
  cnt_to(63 downto 48) <= integer_to_std_logic_vector(cnt_63_48, 16, op_arith);
  cnt_to(47 downto 32) <= integer_to_std_logic_vector(cnt_47_32, 16, op_arith);
  cnt_to(31 downto 16) <= integer_to_std_logic_vector(cnt_31_16, 16, op_arith);
  cnt_to(15 downto 0) <= integer_to_std_logic_vector(cnt_15_0, 16, op_arith);
  op <= op_net;
  core_ce <= ce and en(0);
  rst_overrides_en <= rst(0) or en(0);
  limit : if (count_limited = 1) generate
    eq_cnt_to : process (op_net, cnt_to)
    begin
      op_thresh0 <= equals(op_net, cnt_to(op_width - 1 downto 0),
                     op_width, op_arith);
    end process;
    core_sinit <= (op_thresh0 or clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  no_limit : if (count_limited = 0) generate
    core_sinit <= (clr or rst(0)) and ce and rst_overrides_en;
  end generate;
  comp0: if ((core_name0 = "cntr_11_0_bcc28bfecf25caff")) generate
    core_instance0: cntr_11_0_bcc28bfecf25caff
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_86806e294f737f4c")) generate
    core_instance1: cntr_11_0_86806e294f737f4c
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp2: if ((core_name0 = "cntr_11_0_36e2bb554c95560d")) generate
    core_instance2: cntr_11_0_36e2bb554c95560d
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp3: if ((core_name0 = "cntr_11_0_f068fb73312ae1e5")) generate
    core_instance3: cntr_11_0_f068fb73312ae1e5
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp4: if ((core_name0 = "cntr_11_0_d24951bef2f0cdc9")) generate
    core_instance4: cntr_11_0_d24951bef2f0cdc9
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c5804edea5 is
  port (
    in0 : in std_logic_vector((16 - 1) downto 0);
    in1 : in std_logic_vector((4 - 1) downto 0);
    in2 : in std_logic_vector((9 - 1) downto 0);
    in3 : in std_logic_vector((3 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c5804edea5;


architecture behavior of concat_c5804edea5 is
  signal in0_1_23: unsigned((16 - 1) downto 0);
  signal in1_1_27: unsigned((4 - 1) downto 0);
  signal in2_1_31: unsigned((9 - 1) downto 0);
  signal in3_1_35: unsigned((3 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6293007044 is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6293007044;


architecture behavior of constant_6293007044 is
begin
  op <= "1";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_822933f89b is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_822933f89b;


architecture behavior of constant_822933f89b is
begin
  op <= "000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9f5572ba51 is
  port (
    op : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9f5572ba51;


architecture behavior of constant_9f5572ba51 is
begin
  op <= "0000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c4c603edf2 is
  port (
    op : out std_logic_vector((64 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c4c603edf2;


architecture behavior of constant_c4c603edf2 is
begin
  op <= "0000000000000000000000000000000000000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_91ef1678ca is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_91ef1678ca;


architecture behavior of constant_91ef1678ca is
begin
  op <= "00000000";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_129040d58e is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((5 - 1) downto 0);
    d1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_129040d58e;


architecture behavior of mux_129040d58e is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((5 - 1) downto 0);
  signal d1_1_27: std_logic_vector((9 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((9 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 9, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_82fb466a8b is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_82fb466a8b;


architecture behavior of relational_82fb466a8b is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
entity xlcounter_free_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free_wlan_phy_tx_pmd ;
architecture behavior of xlcounter_free_wlan_phy_tx_pmd is
  component cntr_11_0_36e2bb554c95560d
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_36e2bb554c95560d:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_36e2bb554c95560d:
    component is "true";
  attribute box_type of cntr_11_0_36e2bb554c95560d:
    component  is "black_box";
  component cntr_11_0_6454489cfe866515
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_6454489cfe866515:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_6454489cfe866515:
    component is "true";
  attribute box_type of cntr_11_0_6454489cfe866515:
    component  is "black_box";
  component cntr_11_0_d24951bef2f0cdc9
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d24951bef2f0cdc9:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d24951bef2f0cdc9:
    component is "true";
  attribute box_type of cntr_11_0_d24951bef2f0cdc9:
    component  is "black_box";
  component cntr_11_0_d66925a45384983e
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_d66925a45384983e:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_d66925a45384983e:
    component is "true";
  attribute box_type of cntr_11_0_d66925a45384983e:
    component  is "black_box";
  component cntr_11_0_f068fb73312ae1e5
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_f068fb73312ae1e5:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_f068fb73312ae1e5:
    component is "true";
  attribute box_type of cntr_11_0_f068fb73312ae1e5:
    component  is "black_box";
  component cntr_11_0_86806e294f737f4c
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of cntr_11_0_86806e294f737f4c:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_86806e294f737f4c:
    component is "true";
  attribute box_type of cntr_11_0_86806e294f737f4c:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_36e2bb554c95560d")) generate
    core_instance0: cntr_11_0_36e2bb554c95560d
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp1: if ((core_name0 = "cntr_11_0_6454489cfe866515")) generate
    core_instance1: cntr_11_0_6454489cfe866515
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp2: if ((core_name0 = "cntr_11_0_d24951bef2f0cdc9")) generate
    core_instance2: cntr_11_0_d24951bef2f0cdc9
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp3: if ((core_name0 = "cntr_11_0_d66925a45384983e")) generate
    core_instance3: cntr_11_0_d66925a45384983e
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp4: if ((core_name0 = "cntr_11_0_f068fb73312ae1e5")) generate
    core_instance4: cntr_11_0_f068fb73312ae1e5
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
  comp5: if ((core_name0 = "cntr_11_0_86806e294f737f4c")) generate
    core_instance5: cntr_11_0_86806e294f737f4c
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_b0082e75ff is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    d5 : in std_logic_vector((1 - 1) downto 0);
    d6 : in std_logic_vector((1 - 1) downto 0);
    d7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_b0082e75ff;


architecture behavior of mux_b0082e75ff is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal d3_1_33: std_logic_vector((1 - 1) downto 0);
  signal d4_1_36: std_logic_vector((1 - 1) downto 0);
  signal d5_1_39: std_logic_vector((1 - 1) downto 0);
  signal d6_1_42: std_logic_vector((1 - 1) downto 0);
  signal d7_1_45: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((1 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_c762ea476a is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    d2 : in std_logic_vector((8 - 1) downto 0);
    d3 : in std_logic_vector((8 - 1) downto 0);
    d4 : in std_logic_vector((8 - 1) downto 0);
    d5 : in std_logic_vector((8 - 1) downto 0);
    d6 : in std_logic_vector((8 - 1) downto 0);
    d7 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_c762ea476a;


architecture behavior of mux_c762ea476a is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal d2_1_30: std_logic_vector((8 - 1) downto 0);
  signal d3_1_33: std_logic_vector((8 - 1) downto 0);
  signal d4_1_36: std_logic_vector((8 - 1) downto 0);
  signal d5_1_39: std_logic_vector((8 - 1) downto 0);
  signal d6_1_42: std_logic_vector((8 - 1) downto 0);
  signal d7_1_45: std_logic_vector((8 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((8 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_cda50df78a is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_cda50df78a;


architecture behavior of constant_cda50df78a is
begin
  op <= "00";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1d6ad1c713 is
  port (
    op : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1d6ad1c713;


architecture behavior of constant_1d6ad1c713 is
begin
  op <= "111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_a10351e9f3 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((3 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    d2 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((3 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_a10351e9f3;


architecture behavior of mux_a10351e9f3 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((3 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal d2_1_30: std_logic_vector((2 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((3 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= cast(d1_1_27, 0, 3, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= cast(d2_1_30, 0, 3, 0, xlUnsigned);
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_8fc7f5539b is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_8fc7f5539b;


architecture behavior of relational_8fc7f5539b is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_632978e9ce is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((3 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_632978e9ce;


architecture behavior of relational_632978e9ce is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((3 - 1) downto 0);
  signal cast_12_12: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_12 <= u2u_cast(a_1_31, 0, 3, 0);
  result_12_3_rel <= cast_12_12 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_7673b9b993 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    in4 : in std_logic_vector((1 - 1) downto 0);
    in5 : in std_logic_vector((1 - 1) downto 0);
    in6 : in std_logic_vector((1 - 1) downto 0);
    in7 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_7673b9b993;


architecture behavior of concat_7673b9b993 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal in4_1_39: unsigned((1 - 1) downto 0);
  signal in5_1_43: unsigned((1 - 1) downto 0);
  signal in6_1_47: unsigned((1 - 1) downto 0);
  signal in7_1_51: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  in4_1_39 <= std_logic_vector_to_unsigned(in4);
  in5_1_43 <= std_logic_vector_to_unsigned(in5);
  in6_1_47 <= std_logic_vector_to_unsigned(in6);
  in7_1_51 <= std_logic_vector_to_unsigned(in7);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35) & unsigned_to_std_logic_vector(in4_1_39) & unsigned_to_std_logic_vector(in5_1_43) & unsigned_to_std_logic_vector(in6_1_47) & unsigned_to_std_logic_vector(in7_1_51));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_dist_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    addr_width: integer := 2;
    latency: integer := 0;
    c_width: integer := 12;
    c_address_width: integer := 4
  );
  port (
    addr: in std_logic_vector(addr_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_dist_wlan_phy_tx_pmd ;
architecture behavior of xlsprom_dist_wlan_phy_tx_pmd is
  component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i           : in std_logic_vector(width - 1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width - 1 downto 0));
  end component;
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  constant num_extra_addr_bits: integer := (c_address_width - addr_width);
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_ce: std_logic;
  component dmg_72_134e91999cae8947
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_134e91999cae8947:
    component is true;
  attribute fpga_dont_touch of dmg_72_134e91999cae8947:
    component is "true";
  attribute box_type of dmg_72_134e91999cae8947:
    component  is "black_box";
  component dmg_72_5efcdb43c0011b51
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      spo: out std_logic_vector(c_width - 1 downto 0) 
    );
  end component;

  attribute syn_black_box of dmg_72_5efcdb43c0011b51:
    component is true;
  attribute fpga_dont_touch of dmg_72_5efcdb43c0011b51:
    component is "true";
  attribute box_type of dmg_72_5efcdb43c0011b51:
    component  is "black_box";
  component dmg_72_28ec6cac12d9767d
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_28ec6cac12d9767d:
    component is true;
  attribute fpga_dont_touch of dmg_72_28ec6cac12d9767d:
    component is "true";
  attribute box_type of dmg_72_28ec6cac12d9767d:
    component  is "black_box";
  component dmg_72_140171b6b191950b
    port (
      a: in std_logic_vector(c_address_width - 1 downto 0);
      clk: in std_logic;
      qspo_ce: in std_logic;
      qspo: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of dmg_72_140171b6b191950b:
    component is true;
  attribute fpga_dont_touch of dmg_72_140171b6b191950b:
    component is "true";
  attribute box_type of dmg_72_140171b6b191950b:
    component  is "black_box";
begin
  need_to_pad_addr: if num_extra_addr_bits > 0 generate
      core_addr(c_address_width - 1 downto addr_width) <= (others => '0');
    core_addr(addr_width - 1 downto 0) <= addr;
  end generate;
  no_need_to_pad_addr: if num_extra_addr_bits = 0 generate
    core_addr <= addr;
  end generate;
  core_ce <= ce and en(0);
  comp0: if ((core_name0 = "dmg_72_134e91999cae8947")) generate
    core_instance0: dmg_72_134e91999cae8947
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp1: if ((core_name0 = "dmg_72_5efcdb43c0011b51")) generate
    core_instance1: dmg_72_5efcdb43c0011b51
      port map (
        a => core_addr,
        spo => core_data_out
      );
  end generate;
  comp2: if ((core_name0 = "dmg_72_28ec6cac12d9767d")) generate
    core_instance2: dmg_72_28ec6cac12d9767d
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  comp3: if ((core_name0 = "dmg_72_140171b6b191950b")) generate
    core_instance3: dmg_72_140171b6b191950b
      port map (
        a => core_addr,
        clk => clk,
        qspo_ce => core_ce,
        qspo => core_data_out
      );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_0_or_1: if (latency <= 1)
  generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a1e126f11c is
  port (
    in0 : in std_logic_vector((8 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    in2 : in std_logic_vector((8 - 1) downto 0);
    in3 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a1e126f11c;


architecture behavior of concat_a1e126f11c is
  signal in0_1_23: unsigned((8 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal in2_1_31: unsigned((8 - 1) downto 0);
  signal in3_1_35: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c048fbe4a5 is
  port (
    in0 : in std_logic_vector((24 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c048fbe4a5;


architecture behavior of concat_c048fbe4a5 is
  signal in0_1_23: unsigned((24 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_6a3d3dd4e5 is
  port (
    ip : in std_logic_vector((32 - 1) downto 0);
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_6a3d3dd4e5;


architecture behavior of inverter_6a3d3dd4e5 is
  signal ip_1_26: unsigned((32 - 1) downto 0);
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of unsigned((32 - 1) downto 0);
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => "00000000000000000000000000000000");
  signal op_mem_22_20_front_din: unsigned((32 - 1) downto 0);
  signal op_mem_22_20_back: unsigned((32 - 1) downto 0);
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: unsigned((32 - 1) downto 0);
begin
  ip_1_26 <= std_logic_vector_to_unsigned(ip);
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= std_logic_vector_to_unsigned(not unsigned_to_std_logic_vector(ip_1_26));
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(internal_ip_12_1_bitnot);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_59f8d33339 is
  port (
    d0 : in std_logic_vector((8 - 1) downto 0);
    d1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_59f8d33339;


architecture behavior of logical_59f8d33339 is
  signal d0_1_24: std_logic_vector((8 - 1) downto 0);
  signal d1_1_27: std_logic_vector((8 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((8 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_b23aa74086 is
  port (
    d0 : in std_logic_vector((32 - 1) downto 0);
    d1 : in std_logic_vector((32 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_b23aa74086;


architecture behavior of logical_b23aa74086 is
  signal d0_1_24: std_logic_vector((32 - 1) downto 0);
  signal d1_1_27: std_logic_vector((32 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((32 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_37567836aa is
  port (
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_37567836aa;


architecture behavior of constant_37567836aa is
begin
  op <= "00000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f3924dc817 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((64 - 1) downto 0);
    d1 : in std_logic_vector((32 - 1) downto 0);
    d2 : in std_logic_vector((32 - 1) downto 0);
    y : out std_logic_vector((64 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f3924dc817;


architecture behavior of mux_f3924dc817 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((64 - 1) downto 0);
  signal d1_1_27: std_logic_vector((32 - 1) downto 0);
  signal d2_1_30: std_logic_vector((32 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((64 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= cast(d1_1_27, 0, 64, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= cast(d2_1_30, 0, 64, 0, xlUnsigned);
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a0c7cd7a34 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    in2 : in std_logic_vector((1 - 1) downto 0);
    in3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a0c7cd7a34;


architecture behavior of concat_a0c7cd7a34 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal in2_1_31: unsigned((1 - 1) downto 0);
  signal in3_1_35: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((4 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  in2_1_31 <= std_logic_vector_to_unsigned(in2);
  in3_1_35 <= std_logic_vector_to_unsigned(in3);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27) & unsigned_to_std_logic_vector(in2_1_31) & unsigned_to_std_logic_vector(in3_1_35));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_d6e645765a is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_d6e645765a;


architecture behavior of constant_d6e645765a is
begin
  op <= "011001000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_c49d820dc8 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_c49d820dc8;


architecture behavior of relational_c49d820dc8 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_14_17: unsigned((6 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_14_17 <= u2u_cast(b_1_34, 0, 6, 0);
  result_14_3_rel <= a_1_31 /= cast_14_17;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_43590be5cb is
  port (
    a : in std_logic_vector((12 - 1) downto 0);
    b : in std_logic_vector((12 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_43590be5cb;


architecture behavior of relational_43590be5cb is
  signal a_1_31: unsigned((12 - 1) downto 0);
  signal b_1_34: unsigned((12 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mcode_block_b45edf5eb5 is
  port (
    signal_rate : in std_logic_vector((4 - 1) downto 0);
    mod_order : out std_logic_vector((3 - 1) downto 0);
    code_rate : out std_logic_vector((2 - 1) downto 0);
    n_cbps : out std_logic_vector((9 - 1) downto 0);
    n_dbps : out std_logic_vector((8 - 1) downto 0);
    valid : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mcode_block_b45edf5eb5;


architecture behavior of mcode_block_b45edf5eb5 is
  signal signal_rate_1_80: unsigned((4 - 1) downto 0);
  signal mod_order_join_39_1: unsigned((3 - 1) downto 0);
  signal n_cbps_join_39_1: unsigned((9 - 1) downto 0);
  signal code_rate_join_39_1: unsigned((2 - 1) downto 0);
  signal valid_join_39_1: unsigned((1 - 1) downto 0);
  signal n_dbps_join_39_1: unsigned((8 - 1) downto 0);
begin
  signal_rate_1_80 <= std_logic_vector_to_unsigned(signal_rate);
  proc_switch_39_1: process (signal_rate_1_80)
  is
  begin
    case signal_rate_1_80 is 
      when "1101" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("001");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("000110000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("00");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("00011000");
      when "1111" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("001");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("000110000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("10");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("00100100");
      when "0101" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("010");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("001100000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("00");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("00110000");
      when "0111" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("010");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("001100000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("10");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("01001000");
      when "1001" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("100");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("011000000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("00");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("01100000");
      when "1011" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("100");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("011000000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("10");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("10010000");
      when "0001" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("110");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("100100000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("01");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("11000000");
      when "0011" =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("110");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("100100000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("10");
        valid_join_39_1 <= std_logic_vector_to_unsigned("1");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("11011000");
      when others =>
        mod_order_join_39_1 <= std_logic_vector_to_unsigned("001");
        n_cbps_join_39_1 <= std_logic_vector_to_unsigned("000110000");
        code_rate_join_39_1 <= std_logic_vector_to_unsigned("00");
        valid_join_39_1 <= std_logic_vector_to_unsigned("0");
        n_dbps_join_39_1 <= std_logic_vector_to_unsigned("00011000");
    end case;
  end process proc_switch_39_1;
  mod_order <= unsigned_to_std_logic_vector(mod_order_join_39_1);
  code_rate <= unsigned_to_std_logic_vector(code_rate_join_39_1);
  n_cbps <= unsigned_to_std_logic_vector(n_cbps_join_39_1);
  n_dbps <= unsigned_to_std_logic_vector(n_dbps_join_39_1);
  valid <= unsigned_to_std_logic_vector(valid_join_39_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c936744458 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c936744458;


architecture behavior of constant_c936744458 is
begin
  op <= "01111000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_a6d07705dd is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_a6d07705dd;


architecture behavior of logical_a6d07705dd is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal d3_1_33: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  d3_1_33 <= d3(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27 or d2_1_30 or d3_1_33;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5a9c998b07 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5a9c998b07;


architecture behavior of relational_5a9c998b07 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_19bf67ea71 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_19bf67ea71;


architecture behavior of relational_19bf67ea71 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal cast_12_12: unsigned((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_12 <= u2u_cast(a_1_31, 0, 9, 0);
  result_12_3_rel <= cast_12_12 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_6cb8f0ce02 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_6cb8f0ce02;


architecture behavior of logical_6cb8f0ce02 is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27 or d2_1_30;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity axi_sgiface is
    generic (
        -- AXI specific.
        -- TODO: need to figure out a way to pass these generics from outside
        C_S_AXI_SUPPORT_BURST   : integer := 0;
        -- TODO: fix the internal ID width to 8
        C_S_AXI_ID_WIDTH        : integer := 8;
        C_S_AXI_DATA_WIDTH      : integer := 32;
        C_S_AXI_ADDR_WIDTH      : integer := 32;
        C_S_AXI_TOTAL_ADDR_LEN  : integer := 12;
        C_S_AXI_LINEAR_ADDR_LEN : integer := 8;
        C_S_AXI_BANK_ADDR_LEN   : integer := 2;
        C_S_AXI_AWLEN_WIDTH     : integer := 8;
        C_S_AXI_ARLEN_WIDTH     : integer := 8
    );
    port (
        -- General.
        AXI_AClk      : in  std_logic;
        AXI_AResetN    : in  std_logic;
        -- not used
        AXI_Ce        : in  std_logic;
  
        -- AXI Port.
        S_AXI_AWADDR  : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_AWID    : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_AWLEN   : in  std_logic_vector(C_S_AXI_AWLEN_WIDTH-1 downto 0);
        S_AXI_AWSIZE  : in  std_logic_vector(2 downto 0);
        S_AXI_AWBURST : in  std_logic_vector(1 downto 0);
        S_AXI_AWLOCK  : in  std_logic_vector(1 downto 0);
        S_AXI_AWCACHE : in  std_logic_vector(3 downto 0);
        S_AXI_AWPROT  : in  std_logic_vector(2 downto 0);
        S_AXI_AWVALID : in  std_logic;
        S_AXI_AWREADY : out std_logic;
        
        S_AXI_WLAST   : in  std_logic;
        S_AXI_WDATA   : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_WSTRB   : in  std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
        S_AXI_WVALID  : in  std_logic;
        S_AXI_WREADY  : out std_logic;
        
        S_AXI_BRESP   : out std_logic_vector(1 downto 0);
        S_AXI_BID     : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_BVALID  : out std_logic;
        S_AXI_BREADY  : in  std_logic;
        
        S_AXI_ARADDR  : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_ARID    : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_ARLEN   : in  std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
        S_AXI_ARSIZE  : in  std_logic_vector(2 downto 0);
        S_AXI_ARBURST : in  std_logic_vector(1 downto 0);
        S_AXI_ARLOCK  : in  std_logic_vector(1 downto 0);
        S_AXI_ARCACHE : in  std_logic_vector(3 downto 0);
        S_AXI_ARPROT  : in  std_logic_vector(2 downto 0);
        S_AXI_ARVALID : in  std_logic;
        S_AXI_ARREADY : out std_logic;
        
        -- 'From Register'
        -- 'STATUS'
        sm_STATUS_dout : in std_logic_vector(32-1 downto 0);
        -- 'To Register'
        -- 'Timing'
        sm_Timing_dout : in std_logic_vector(32-1 downto 0);
        sm_Timing_din  : out std_logic_vector(32-1 downto 0);
        sm_Timing_en   : out std_logic;
        -- 'Config'
        sm_Config_dout : in std_logic_vector(32-1 downto 0);
        sm_Config_din  : out std_logic_vector(32-1 downto 0);
        sm_Config_en   : out std_logic;
        -- 'PKT_BUF_SEL'
        sm_PKT_BUF_SEL_dout : in std_logic_vector(32-1 downto 0);
        sm_PKT_BUF_SEL_din  : out std_logic_vector(32-1 downto 0);
        sm_PKT_BUF_SEL_en   : out std_logic;
        -- 'Output_Scaling'
        sm_Output_Scaling_dout : in std_logic_vector(32-1 downto 0);
        sm_Output_Scaling_din  : out std_logic_vector(32-1 downto 0);
        sm_Output_Scaling_en   : out std_logic;
        -- 'TX_START'
        sm_TX_START_dout : in std_logic_vector(32-1 downto 0);
        sm_TX_START_din  : out std_logic_vector(32-1 downto 0);
        sm_TX_START_en   : out std_logic;
        -- 'FFT_Config'
        sm_FFT_Config_dout : in std_logic_vector(32-1 downto 0);
        sm_FFT_Config_din  : out std_logic_vector(32-1 downto 0);
        sm_FFT_Config_en   : out std_logic;
        -- 'From FIFO'
        -- 'To FIFO'
        -- 'Shared Memory'

        S_AXI_RLAST   : out std_logic;
        S_AXI_RID     : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
        S_AXI_RDATA   : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_RRESP   : out std_logic_vector(1 downto 0);
        S_AXI_RVALID  : out std_logic;
        S_AXI_RREADY  : in  std_logic
    );
end entity axi_sgiface;

architecture IMP of axi_sgiface is

-- Internal signals for write channel.
signal S_AXI_BVALID_i       : std_logic;
signal S_AXI_BID_i          : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
signal S_AXI_WREADY_i       : std_logic;
  
-- Internal signals for read channels.
signal S_AXI_ARLEN_i        : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
signal S_AXI_RLAST_i        : std_logic;
signal S_AXI_RREADY_i       : std_logic;
signal S_AXI_RVALID_i       : std_logic;
signal S_AXI_RDATA_i        : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal S_AXI_RID_i          : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);

-- for read channel
signal read_bank_addr_i     : std_logic_vector(C_S_AXI_BANK_ADDR_LEN-1 downto 0);
signal read_linear_addr_i   : std_logic_vector(C_S_AXI_LINEAR_ADDR_LEN-1 downto 0);
-- for write channel
signal write_bank_addr_i    : std_logic_vector(C_S_AXI_BANK_ADDR_LEN-1 downto 0);
signal write_linear_addr_i  : std_logic_vector(C_S_AXI_LINEAR_ADDR_LEN-1 downto 0);

signal reg_bank_out_i       : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal fifo_bank_out_i      : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal shmem_bank_out_i     : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
    
-- 'From Register'
-- 'STATUS'
signal sm_STATUS_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'To Register'
-- 'Timing'
signal sm_Timing_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Timing_en_i    : std_logic;
signal sm_Timing_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'Config'
signal sm_Config_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Config_en_i    : std_logic;
signal sm_Config_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'PKT_BUF_SEL'
signal sm_PKT_BUF_SEL_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_PKT_BUF_SEL_en_i    : std_logic;
signal sm_PKT_BUF_SEL_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'Output_Scaling'
signal sm_Output_Scaling_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_Output_Scaling_en_i    : std_logic;
signal sm_Output_Scaling_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'TX_START'
signal sm_TX_START_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_TX_START_en_i    : std_logic;
signal sm_TX_START_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'FFT_Config'
signal sm_FFT_Config_din_i   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
signal sm_FFT_Config_en_i    : std_logic;
signal sm_FFT_Config_dout_i  : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
-- 'From FIFO'
-- 'To FIFO'
-- 'Shared Memory'

type t_read_state is (IDLE, READ_PREP, READ_DATA);
signal read_state : t_read_state;

type t_write_state is (IDLE, WRITE_DATA, WRITE_RESPONSE);
signal write_state : t_write_state;

type t_memmap_state is (READ, WRITE);
signal memmap_state : t_memmap_state;

constant C_READ_PREP_DELAY : std_logic_vector(1 downto 0) := "11";

signal read_prep_counter : std_logic_vector(1 downto 0);
signal read_addr_counter : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);
signal read_data_counter : std_logic_vector(C_S_AXI_ARLEN_WIDTH-1 downto 0);

-- enable of shared BRAMs
signal s_shram_en : std_logic;

signal write_addr_valid : std_logic;
signal write_ready : std_logic;

-- 're' of From/To FIFOs
signal s_fifo_re : std_logic;
-- 'we' of To FIFOs
signal s_fifo_we : std_logic;

begin

-- enable for 'Shared Memory' blocks

-- conversion to match with the data bus width
-- 'From Register'
-- 'STATUS'
gen_sm_STATUS_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_STATUS_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_STATUS_dout_i;
sm_STATUS_dout_i(32-1 downto 0) <= sm_STATUS_dout;
-- 'To Register'
-- 'Timing'
sm_Timing_din     <= sm_Timing_din_i(32-1 downto 0);
sm_Timing_en      <= sm_Timing_en_i;
gen_sm_Timing_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Timing_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Timing_dout_i;
sm_Timing_dout_i(32-1 downto 0) <= sm_Timing_dout;
-- 'Config'
sm_Config_din     <= sm_Config_din_i(32-1 downto 0);
sm_Config_en      <= sm_Config_en_i;
gen_sm_Config_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Config_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Config_dout_i;
sm_Config_dout_i(32-1 downto 0) <= sm_Config_dout;
-- 'PKT_BUF_SEL'
sm_PKT_BUF_SEL_din     <= sm_PKT_BUF_SEL_din_i(32-1 downto 0);
sm_PKT_BUF_SEL_en      <= sm_PKT_BUF_SEL_en_i;
gen_sm_PKT_BUF_SEL_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_PKT_BUF_SEL_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_PKT_BUF_SEL_dout_i;
sm_PKT_BUF_SEL_dout_i(32-1 downto 0) <= sm_PKT_BUF_SEL_dout;
-- 'Output_Scaling'
sm_Output_Scaling_din     <= sm_Output_Scaling_din_i(32-1 downto 0);
sm_Output_Scaling_en      <= sm_Output_Scaling_en_i;
gen_sm_Output_Scaling_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_Output_Scaling_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_Output_Scaling_dout_i;
sm_Output_Scaling_dout_i(32-1 downto 0) <= sm_Output_Scaling_dout;
-- 'TX_START'
sm_TX_START_din     <= sm_TX_START_din_i(32-1 downto 0);
sm_TX_START_en      <= sm_TX_START_en_i;
gen_sm_TX_START_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_TX_START_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_TX_START_dout_i;
sm_TX_START_dout_i(32-1 downto 0) <= sm_TX_START_dout;
-- 'FFT_Config'
sm_FFT_Config_din     <= sm_FFT_Config_din_i(32-1 downto 0);
sm_FFT_Config_en      <= sm_FFT_Config_en_i;
gen_sm_FFT_Config_dout_i: if (32 < C_S_AXI_DATA_WIDTH) generate
    sm_FFT_Config_dout_i(C_S_AXI_DATA_WIDTH-1 downto 32) <= (others => '0');
end generate gen_sm_FFT_Config_dout_i;
sm_FFT_Config_dout_i(32-1 downto 0) <= sm_FFT_Config_dout;
-- 'From FIFO'
-- 'To FIFO'
-- 'Shared Memory'

ReadWriteSelect: process(memmap_state) is begin
    if (memmap_state = READ) then
    else
    end if;
end process ReadWriteSelect;

-----------------------------------------------------------------------------
-- address for 'Shared Memory'
-----------------------------------------------------------------------------
SharedMemory_Addr_ResetN : process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            memmap_state <= READ;
        else
            if (S_AXI_AWVALID = '1') then
                -- write operation
                memmap_state <= WRITE;
            elsif (S_AXI_ARVALID = '1') then
                -- read operation
                memmap_state <= READ;
            end if;
        end if;
    end if;
end process SharedMemory_Addr_ResetN;

-----------------------------------------------------------------------------
-- WRITE Command Control
-----------------------------------------------------------------------------
S_AXI_BID     <= S_AXI_BID_i;
S_AXI_BVALID  <= S_AXI_BVALID_i;
S_AXI_WREADY  <= S_AXI_WREADY_i;
-- No error checking
S_AXI_BRESP  <= (others=>'0');

PROC_AWREADY_ACK: process(read_state, write_state, S_AXI_ARVALID, S_AXI_AWVALID) is begin
    if (write_state = IDLE and S_AXI_AWVALID = '1' and read_state = IDLE) then
        S_AXI_AWREADY <= S_AXI_AWVALID;
    else
        S_AXI_AWREADY <= '0';
    end if;
end process PROC_AWREADY_ACK;

Cmd_Decode_Write: process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            write_addr_valid    <= '0';
            write_ready         <= '0';
            s_fifo_we           <= '0';
            S_AXI_BVALID_i      <= '0';
            S_AXI_BID_i         <= (others => '0');
            write_bank_addr_i   <= (others => '0');
            write_linear_addr_i <= (others => '0');
        else
            if (write_state = IDLE) then
                if (S_AXI_AWVALID = '1' and read_state = IDLE) then
                    -- reflect awid
                    S_AXI_BID_i <= S_AXI_AWID;

                    -- latch bank and linear addresses
                    write_bank_addr_i   <= S_AXI_AWADDR(C_S_AXI_TOTAL_ADDR_LEN-1 downto C_S_AXI_LINEAR_ADDR_LEN+2);
                    write_linear_addr_i <= S_AXI_AWADDR(C_S_AXI_LINEAR_ADDR_LEN+1 downto 2);
                    write_addr_valid <= '1';
                    s_fifo_we <= '1';

                    -- write state transition
                    write_state <= WRITE_DATA;
                end if;
            elsif (write_state = WRITE_DATA) then
                write_ready <= '1';
                s_fifo_we <= '0';
                write_addr_valid <= S_AXI_WVALID;
                
                if (S_AXI_WVALID = '1' and write_ready = '1') then
                    write_linear_addr_i <= Std_Logic_Vector(unsigned(write_linear_addr_i) + 1);
                end if;

                if (S_AXI_WLAST = '1' and write_ready = '1') then
                    -- start responding through B channel upon the last write data sample
                    S_AXI_BVALID_i <= '1';
                    -- write data is over
                    write_addr_valid <= '0';
                    write_ready <= '0';
                    -- write state transition
                    write_state <= WRITE_RESPONSE;
                end if;
            elsif (write_state = WRITE_RESPONSE) then

                if (S_AXI_BREADY = '1') then
                    -- write respond is over
                    S_AXI_BVALID_i <= '0';
                    S_AXI_BID_i <= (others => '0');

                    -- write state transition
                    write_state <= IDLE;
                end if;
            end if;
        end if;
    end if;
end process Cmd_Decode_Write;

Write_Linear_Addr_Decode : process(AXI_AClk) is 

begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            -- 'To Register'
            -- Timing din/en
            sm_Timing_din_i <= (others => '0');
            sm_Timing_en_i <= '0';
            -- Config din/en
            sm_Config_din_i <= (others => '0');
            sm_Config_en_i <= '0';
            -- PKT_BUF_SEL din/en
            sm_PKT_BUF_SEL_din_i <= (others => '0');
            sm_PKT_BUF_SEL_en_i <= '0';
            -- Output_Scaling din/en
            sm_Output_Scaling_din_i <= (others => '0');
            sm_Output_Scaling_en_i <= '0';
            -- TX_START din/en
            sm_TX_START_din_i <= (others => '0');
            sm_TX_START_en_i <= '0';
            -- FFT_Config din/en
            sm_FFT_Config_din_i <= (others => '0');
            sm_FFT_Config_en_i <= '0';
            -- 'To FIFO'
            -- 'Shared Memory'
        else
            -- default assignments

            -- 'To Register'
            if (unsigned(write_bank_addr_i) = 2) then
                if (unsigned(write_linear_addr_i) = 0) then
                    -- Timing din/en
                    sm_Timing_din_i <= S_AXI_WDATA;
                    sm_Timing_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 1) then
                    -- Config din/en
                    sm_Config_din_i <= S_AXI_WDATA;
                    sm_Config_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 2) then
                    -- PKT_BUF_SEL din/en
                    sm_PKT_BUF_SEL_din_i <= S_AXI_WDATA;
                    sm_PKT_BUF_SEL_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 3) then
                    -- Output_Scaling din/en
                    sm_Output_Scaling_din_i <= S_AXI_WDATA;
                    sm_Output_Scaling_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 4) then
                    -- TX_START din/en
                    sm_TX_START_din_i <= S_AXI_WDATA;
                    sm_TX_START_en_i  <= write_addr_valid;
                elsif (unsigned(write_linear_addr_i) = 5) then
                    -- FFT_Config din/en
                    sm_FFT_Config_din_i <= S_AXI_WDATA;
                    sm_FFT_Config_en_i  <= write_addr_valid;
                end if;
            end if;        
        
        
        end if;
    end if;
end process Write_Linear_Addr_Decode;
 
-----------------------------------------------------------------------------
-- READ Control
-----------------------------------------------------------------------------

S_AXI_RDATA  <= S_AXI_RDATA_i;
S_AXI_RVALID  <= S_AXI_RVALID_i;
S_AXI_RLAST   <= S_AXI_RLAST_i;
S_AXI_RID     <= S_AXI_RID_i;
-- TODO: no error checking
S_AXI_RRESP <= (others=>'0');

PROC_ARREADY_ACK: process(read_state, S_AXI_ARVALID, write_state, S_AXI_AWVALID) is begin
    -- Note: WRITE has higher priority than READ
    if (read_state = IDLE and S_AXI_ARVALID = '1' and write_state = IDLE and S_AXI_AWVALID /= '1') then
        S_AXI_ARREADY <= S_AXI_ARVALID;
    else
        S_AXI_ARREADY <= '0';
    end if;
end process PROC_ARREADY_ACK;

S_AXI_WREADY_i <= write_ready;

Process_Sideband: process(write_state, read_state) is begin
    if (read_state = READ_PREP) then
        s_shram_en <= '1';
    elsif (read_state = READ_DATA) then
        s_shram_en <= S_AXI_RREADY;
    elsif (write_state = WRITE_DATA) then
        s_shram_en <= S_AXI_WVALID;
    else
        s_shram_en <= '0';
    end if;
end process Process_Sideband;

Cmd_Decode_Read: process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            S_AXI_RVALID_i <= '0';
            read_bank_addr_i    <= (others => '0');
            read_linear_addr_i  <= (others => '0');
            S_AXI_ARLEN_i       <= (others => '0');
            S_AXI_RLAST_i       <= '0';
            S_AXI_RID_i         <= (others => '0');
            read_state          <= IDLE;
            read_prep_counter   <= (others => '0');
            read_addr_counter   <= (others => '0');
            read_data_counter   <= (others => '0');
        else
            -- default assignments
            s_fifo_re <= '0';

            if (read_state = IDLE) then
                -- Note WRITE has higher priority than READ
                if (S_AXI_ARVALID = '1' and write_state = IDLE and S_AXI_AWVALID /= '1') then
                    -- extract bank and linear addresses
                    read_bank_addr_i    <= S_AXI_ARADDR(C_S_AXI_TOTAL_ADDR_LEN-1 downto C_S_AXI_LINEAR_ADDR_LEN+2);
                    read_linear_addr_i  <= S_AXI_ARADDR(C_S_AXI_LINEAR_ADDR_LEN+1 downto 2);
                    s_fifo_re <= '1';

                    -- reflect arid
                    S_AXI_RID_i <= S_AXI_ARID;

                    -- load read liner address and data counter
                    read_addr_counter <= S_AXI_ARLEN;
                    read_data_counter <= S_AXI_ARLEN;

                    -- load read preparation counter
                    read_prep_counter <= C_READ_PREP_DELAY;
                    -- read state transition
                    read_state <= READ_PREP;
                end if;
            elsif (read_state = READ_PREP) then
                if (unsigned(read_prep_counter) = 0) then
                    if (unsigned(read_data_counter) = 0) then
                        -- tag the last data generated by the slave
                        S_AXI_RLAST_i <= '1';
                    end if;
                    -- valid data appears
                    S_AXI_RVALID_i <= '1';
                    -- read state transition
                    read_state <= READ_DATA;
                else
                    -- decrease read preparation counter
                    read_prep_counter <= Std_Logic_Vector(unsigned(read_prep_counter) - 1);
                end if;

                if (unsigned(read_prep_counter) /= 3 and unsigned(read_addr_counter) /= 0) then
                    -- decrease address counter
                    read_addr_counter <= Std_Logic_Vector(unsigned(read_addr_counter) - 1);
                    -- increase linear address (no band crossing)
                    read_linear_addr_i <= Std_Logic_Vector(unsigned(read_linear_addr_i) + 1);
                end if;
            elsif (read_state = READ_DATA) then
                if (S_AXI_RREADY = '1') then
                    if (unsigned(read_data_counter) = 1) then
                        -- tag the last data generated by the slave
                        S_AXI_RLAST_i <= '1';
                    end if;

                    if (unsigned(read_data_counter) = 0) then
                        -- arid
                        S_AXI_RID_i <= (others => '0');
                        -- rlast
                        S_AXI_RLAST_i <= '0';
                        -- no more valid data
                        S_AXI_RVALID_i <= '0';
                        -- read state transition
                        read_state <= IDLE;
                    else
                        -- decrease read preparation counter
                        read_data_counter <= Std_Logic_Vector(unsigned(read_data_counter) - 1);

                        if (unsigned(read_addr_counter) /= 0) then
                            -- decrease address counter
                            read_addr_counter <= Std_Logic_Vector(unsigned(read_addr_counter) - 1);
                            -- increase linear address (no band crossing)
                            read_linear_addr_i <= Std_Logic_Vector(unsigned(read_linear_addr_i) + 1);
                        end if;
                    end if;
                end if;
            end if;

        end if;
    end if;
end process Cmd_Decode_Read;

Read_Linear_Addr_Decode : process(AXI_AClk) is begin
    if (AXI_AClk'event and AXI_AClk = '1') then
        if (AXI_AResetN = '0') then
            reg_bank_out_i   <= (others => '0');
            fifo_bank_out_i  <= (others => '0');
            shmem_bank_out_i <= (others => '0');
            S_AXI_RDATA_i    <= (others => '0');
        else
            if (unsigned(read_bank_addr_i) = 2) then
                -- 'From Register'
                if (unsigned(read_linear_addr_i) = 6) then
                    -- 'STATUS' dout
                    reg_bank_out_i <= sm_STATUS_dout_i;
                end if;
                -- 'To Register' (with register readback)
                if (unsigned(read_linear_addr_i) = 0) then
                    -- 'Timing' dout
                    reg_bank_out_i <= sm_Timing_dout_i;
                elsif (unsigned(read_linear_addr_i) = 1) then
                    -- 'Config' dout
                    reg_bank_out_i <= sm_Config_dout_i;
                elsif (unsigned(read_linear_addr_i) = 2) then
                    -- 'PKT_BUF_SEL' dout
                    reg_bank_out_i <= sm_PKT_BUF_SEL_dout_i;
                elsif (unsigned(read_linear_addr_i) = 3) then
                    -- 'Output_Scaling' dout
                    reg_bank_out_i <= sm_Output_Scaling_dout_i;
                elsif (unsigned(read_linear_addr_i) = 4) then
                    -- 'TX_START' dout
                    reg_bank_out_i <= sm_TX_START_dout_i;
                elsif (unsigned(read_linear_addr_i) = 5) then
                    -- 'FFT_Config' dout
                    reg_bank_out_i <= sm_FFT_Config_dout_i;
                end if;

                S_AXI_RDATA_i <= reg_bank_out_i;
            elsif (unsigned(read_bank_addr_i) = 1) then
                -- 'From FIFO'
                -- 'To FIFO'

                S_AXI_RDATA_i <= fifo_bank_out_i;
            elsif (unsigned(read_bank_addr_i) = 0 and s_shram_en = '1') then
                -- 'Shared Memory'

                S_AXI_RDATA_i <= shmem_bank_out_i;
            end if;
        end if;
    end if;
end process Read_Linear_Addr_Decode;

end architecture IMP;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity xlfast_fourier_transform_66965782653510ded5a0002b36532651 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    event_data_in_channel_halt:out std_logic;
    event_data_out_channel_halt:out std_logic;
    event_fft_overflow:out std_logic;
    event_frame_started:out std_logic;
    event_status_channel_halt:out std_logic;
    event_tlast_missing:out std_logic;
    event_tlast_unexpected:out std_logic;
    m_axis_data_tdata_xk_im:out std_logic_vector(15 downto 0);
    m_axis_data_tdata_xk_re:out std_logic_vector(15 downto 0);
    m_axis_data_tlast:out std_logic;
    m_axis_data_tready:in std_logic;
    m_axis_data_tuser_ovflo:out std_logic_vector(0 downto 0);
    m_axis_data_tuser_xk_index:out std_logic_vector(5 downto 0);
    m_axis_data_tvalid:out std_logic;
    m_axis_status_tdata_ovflo:out std_logic_vector(0 downto 0);
    m_axis_status_tready:in std_logic;
    m_axis_status_tvalid:out std_logic;
    rst:in std_logic;
    s_axis_config_tdata_cp_len:in std_logic_vector(5 downto 0);
    s_axis_config_tdata_fwd_inv:in std_logic_vector(0 downto 0);
    s_axis_config_tdata_scale_sch:in std_logic_vector(5 downto 0);
    s_axis_config_tready:out std_logic;
    s_axis_config_tvalid:in std_logic;
    s_axis_data_tdata_xn_im:in std_logic_vector(15 downto 0);
    s_axis_data_tdata_xn_re:in std_logic_vector(15 downto 0);
    s_axis_data_tlast:in std_logic;
    s_axis_data_tready:out std_logic;
    s_axis_data_tvalid:in std_logic
  );
end xlfast_fourier_transform_66965782653510ded5a0002b36532651;


architecture behavior of xlfast_fourier_transform_66965782653510ded5a0002b36532651  is
  component xfft_v8_0_6e4d6522fcd78ca0
    port(
      aclk:in std_logic;
      aclken:in std_logic;
      aresetn:in std_logic;
      event_data_in_channel_halt:out std_logic;
      event_data_out_channel_halt:out std_logic;
      event_fft_overflow:out std_logic;
      event_frame_started:out std_logic;
      event_status_channel_halt:out std_logic;
      event_tlast_missing:out std_logic;
      event_tlast_unexpected:out std_logic;
      m_axis_data_tdata:out std_logic_vector(31 downto 0);
      m_axis_data_tlast:out std_logic;
      m_axis_data_tready:in std_logic;
      m_axis_data_tuser:out std_logic_vector(15 downto 0);
      m_axis_data_tvalid:out std_logic;
      m_axis_status_tdata:out std_logic_vector(7 downto 0);
      m_axis_status_tready:in std_logic;
      m_axis_status_tvalid:out std_logic;
      s_axis_config_tdata:in std_logic_vector(15 downto 0);
      s_axis_config_tready:out std_logic;
      s_axis_config_tvalid:in std_logic;
      s_axis_data_tdata:in std_logic_vector(31 downto 0);
      s_axis_data_tlast:in std_logic;
      s_axis_data_tready:out std_logic;
      s_axis_data_tvalid:in std_logic
    );
end component;
signal aresetn_net: std_logic := '0';
signal m_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
signal m_axis_data_tuser_net: std_logic_vector(15 downto 0) := (others=>'0');
signal m_axis_status_tdata_net: std_logic_vector(7 downto 0) := (others=>'0');
signal s_axis_config_tdata_net: std_logic_vector(15 downto 0) := (others=>'0');
signal s_axis_data_tdata_net: std_logic_vector(31 downto 0) := (others=>'0');
begin
  aresetn_net <= rst or (not ce);
  m_axis_data_tdata_xk_im <= m_axis_data_tdata_net(31 downto 16);
  m_axis_data_tdata_xk_re <= m_axis_data_tdata_net(15 downto 0);
  m_axis_data_tuser_ovflo <= m_axis_data_tuser_net(8 downto 8);
  m_axis_data_tuser_xk_index <= m_axis_data_tuser_net(5 downto 0);
  m_axis_status_tdata_ovflo <= m_axis_status_tdata_net(0 downto 0);
  s_axis_config_tdata_net(14 downto 9) <= s_axis_config_tdata_scale_sch;
  s_axis_config_tdata_net(8 downto 8) <= s_axis_config_tdata_fwd_inv;
  s_axis_config_tdata_net(5 downto 0) <= s_axis_config_tdata_cp_len;
  s_axis_data_tdata_net(31 downto 16) <= s_axis_data_tdata_xn_im;
  s_axis_data_tdata_net(15 downto 0) <= s_axis_data_tdata_xn_re;
  xfft_v8_0_6e4d6522fcd78ca0_instance : xfft_v8_0_6e4d6522fcd78ca0
    port map(
      aclk=>clk,
      aclken=>ce,
      aresetn=>aresetn_net,
      event_data_in_channel_halt=>event_data_in_channel_halt,
      event_data_out_channel_halt=>event_data_out_channel_halt,
      event_fft_overflow=>event_fft_overflow,
      event_frame_started=>event_frame_started,
      event_status_channel_halt=>event_status_channel_halt,
      event_tlast_missing=>event_tlast_missing,
      event_tlast_unexpected=>event_tlast_unexpected,
      m_axis_data_tdata=>m_axis_data_tdata_net,
      m_axis_data_tlast=>m_axis_data_tlast,
      m_axis_data_tready=>m_axis_data_tready,
      m_axis_data_tuser=>m_axis_data_tuser_net,
      m_axis_data_tvalid=>m_axis_data_tvalid,
      m_axis_status_tdata=>m_axis_status_tdata_net,
      m_axis_status_tready=>m_axis_status_tready,
      m_axis_status_tvalid=>m_axis_status_tvalid,
      s_axis_config_tdata=>s_axis_config_tdata_net,
      s_axis_config_tready=>s_axis_config_tready,
      s_axis_config_tvalid=>s_axis_config_tvalid,
      s_axis_data_tdata=>s_axis_data_tdata_net,
      s_axis_data_tlast=>s_axis_data_tlast,
      s_axis_data_tready=>s_axis_data_tready,
      s_axis_data_tvalid=>s_axis_data_tvalid
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_a369e00c6b is
  port (
    in0 : in std_logic_vector((16 - 1) downto 0);
    in1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_a369e00c6b;


architecture behavior of concat_a369e00c6b is
  signal in0_1_23: unsigned((16 - 1) downto 0);
  signal in1_1_27: unsigned((16 - 1) downto 0);
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_7025463ea8 is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_7025463ea8;


architecture behavior of reinterpret_7025463ea8 is
  signal input_port_1_40: signed((16 - 1) downto 0);
  signal output_port_5_5_force: unsigned((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_signed(input_port);
  output_port_5_5_force <= signed_to_unsigned(input_port_1_40);
  output_port <= unsigned_to_std_logic_vector(output_port_5_5_force);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_151459306d is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_151459306d;


architecture behavior of reinterpret_151459306d is
  signal input_port_1_40: unsigned((16 - 1) downto 0);
  signal output_port_5_5_force: signed((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port_5_5_force <= unsigned_to_signed(input_port_1_40);
  output_port <= signed_to_std_logic_vector(output_port_5_5_force);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.conv_pkg.all;
entity xlaxififogen_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    tdata_width: integer := -1;
    tdest_width: integer := -1;
    tstrb_width: integer := -1;
    tkeep_width: integer := -1;
    tid_width: integer := -1;
    tuser_width: integer := -1;
    has_aresetn: integer := -1;
    depth_bits: integer :=-1
  );
  port (
      s_aclk: in std_logic;
      ce: in std_logic;
      aresetn: in std_logic;
s_axis_tdata: in std_logic_vector(tdata_width - 1 downto 0):= (others => '0');
s_axis_tdest: in std_logic_vector(tdest_width - 1 downto 0):= (others => '0');
s_axis_tstrb: in std_logic_vector(tstrb_width - 1 downto 0):= (others => '0');
s_axis_tkeep: in std_logic_vector(tkeep_width - 1 downto 0):= (others => '0');
s_axis_tlast: in std_logic := '0';
s_axis_tid  : in std_logic_vector(tid_width - 1 downto 0):= (others => '0');
s_axis_tuser: in std_logic_vector(tuser_width - 1 downto 0):= (others => '0');
m_axis_tdata: out std_logic_vector(tdata_width - 1 downto 0);
m_axis_tdest: out std_logic_vector(tdest_width - 1 downto 0);
m_axis_tstrb: out std_logic_vector(tstrb_width - 1 downto 0);
m_axis_tkeep: out std_logic_vector(tkeep_width - 1 downto 0);
m_axis_tlast: out std_logic;
m_axis_tid  : out std_logic_vector(tid_width - 1 downto 0);
m_axis_tuser: out std_logic_vector(tuser_width - 1 downto 0);
      axis_underflow: out std_logic;
      axis_overflow: out std_logic;
      axis_data_count: out std_logic_vector( depth_bits - 1 downto 0);
      axis_prog_full_thresh: in std_logic_vector( depth_bits - 2 downto 0):= (others => '0');
      axis_prog_empty_thresh: in std_logic_vector(depth_bits - 2 downto 0):= (others => '0');

      s_axis_tvalid: in std_logic;
      s_axis_tready: out std_logic;
      m_axis_tready: in std_logic;
      m_axis_tvalid: out std_logic
  );
end xlaxififogen_wlan_phy_tx_pmd;
architecture behavior of xlaxififogen_wlan_phy_tx_pmd is
  component axififo_fg92_4d50ffea04713b7c
    port (
      s_aclk: in std_logic;
      s_aresetn: in std_logic;
      s_axis_tdata: in std_logic_vector(tdata_width - 1 downto 0);
      s_axis_tlast: in std_logic;
      s_axis_tuser: in std_logic_vector(tuser_width - 1 downto 0);
      s_axis_tvalid: in std_logic;
      s_axis_tready: out std_logic;
      m_axis_tdata: out std_logic_vector(tdata_width - 1 downto 0);
      m_axis_tlast: out std_logic;
      m_axis_tuser: out std_logic_vector(tuser_width - 1 downto 0);
      m_axis_tvalid: out std_logic;
      m_axis_tready: in std_logic

    );
  end component;

  attribute syn_black_box of axififo_fg92_4d50ffea04713b7c:
    component is true;
  attribute fpga_dont_touch of axififo_fg92_4d50ffea04713b7c:
    component is "true";
  attribute box_type of axififo_fg92_4d50ffea04713b7c:
    component  is "black_box";
  signal srst: std_logic:= '0';
  signal reset_gen1: std_logic  := '0';
  signal reset_gen_d1: std_logic        := '0';
  signal reset_gen_d2: std_logic := '0';
begin
  comp0: if ((core_name0 = "axififo_fg92_4d50ffea04713b7c")) generate
    core_instance0: axififo_fg92_4d50ffea04713b7c
      port map (
        s_aclk => s_aclk,
        s_aresetn => srst,
        s_axis_tdata => s_axis_tdata,
        s_axis_tlast => s_axis_tlast,
        s_axis_tuser => s_axis_tuser,
        s_axis_tvalid => s_axis_tvalid,
        s_axis_tready => s_axis_tready,
        m_axis_tdata => m_axis_tdata,
        m_axis_tlast => m_axis_tlast,
        m_axis_tuser => m_axis_tuser,
        m_axis_tvalid => m_axis_tvalid,
        m_axis_tready => m_axis_tready

      );
  end generate;
        srst <= reset_gen_d2 when (has_aresetn = 0)
                else not ( (not aresetn) and ce );
 process(s_aclk)
 begin
         if(s_aclk'event AND s_aclk = '1') then
                         reset_gen1 <= '1';
                         reset_gen_d1 <= reset_gen1;
                         reset_gen_d2 <= reset_gen_d1;
        end if;
 end process;

end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity inverter_e2b989a05e is
  port (
    ip : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end inverter_e2b989a05e;


architecture behavior of inverter_e2b989a05e is
  signal ip_1_26: unsigned((1 - 1) downto 0);
  type array_type_op_mem_22_20 is array (0 to (1 - 1)) of unsigned((1 - 1) downto 0);
  signal op_mem_22_20: array_type_op_mem_22_20 := (
    0 => "0");
  signal op_mem_22_20_front_din: unsigned((1 - 1) downto 0);
  signal op_mem_22_20_back: unsigned((1 - 1) downto 0);
  signal op_mem_22_20_push_front_pop_back_en: std_logic;
  signal internal_ip_12_1_bitnot: unsigned((1 - 1) downto 0);
begin
  ip_1_26 <= std_logic_vector_to_unsigned(ip);
  op_mem_22_20_back <= op_mem_22_20(0);
  proc_op_mem_22_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_22_20_push_front_pop_back_en = '1')) then
        op_mem_22_20(0) <= op_mem_22_20_front_din;
      end if;
    end if;
  end process proc_op_mem_22_20;
  internal_ip_12_1_bitnot <= std_logic_vector_to_unsigned(not unsigned_to_std_logic_vector(ip_1_26));
  op_mem_22_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(internal_ip_12_1_bitnot);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlsprom_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    c_width: integer := 12;
    c_address_width: integer := 4;
    latency: integer := 1
  );
  port (
    addr: in std_logic_vector(c_address_width - 1 downto 0);
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0);
    ce: in std_logic;
    clk: in std_logic;
    data: out std_logic_vector(c_width - 1 downto 0)
  );
end xlsprom_wlan_phy_tx_pmd ;
architecture behavior of xlsprom_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal core_addr: std_logic_vector(c_address_width - 1 downto 0);
  signal core_data_out: std_logic_vector(c_width - 1 downto 0);
  signal core_ce, sinit: std_logic;
  component bmg_72_28f68c2bb9b4d938
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_28f68c2bb9b4d938:
    component is true;
  attribute fpga_dont_touch of bmg_72_28f68c2bb9b4d938:
    component is "true";
  attribute box_type of bmg_72_28f68c2bb9b4d938:
    component  is "black_box";
  component bmg_72_324b883165919716
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_324b883165919716:
    component is true;
  attribute fpga_dont_touch of bmg_72_324b883165919716:
    component is "true";
  attribute box_type of bmg_72_324b883165919716:
    component  is "black_box";
  component bmg_72_f580ae3be5511d30
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_f580ae3be5511d30:
    component is true;
  attribute fpga_dont_touch of bmg_72_f580ae3be5511d30:
    component is "true";
  attribute box_type of bmg_72_f580ae3be5511d30:
    component  is "black_box";
  component bmg_72_3628803596b5ca22
    port (
                              addra: in std_logic_vector(c_address_width - 1 downto 0);
      clka: in std_logic;
      ena: in std_logic;
      douta: out std_logic_vector(c_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of bmg_72_3628803596b5ca22:
    component is true;
  attribute fpga_dont_touch of bmg_72_3628803596b5ca22:
    component is "true";
  attribute box_type of bmg_72_3628803596b5ca22:
    component  is "black_box";
begin
  core_addr <= addr;
  core_ce <= ce and en(0);
  sinit <= rst(0) and ce;
  comp0: if ((core_name0 = "bmg_72_28f68c2bb9b4d938")) generate
    core_instance0: bmg_72_28f68c2bb9b4d938
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp1: if ((core_name0 = "bmg_72_324b883165919716")) generate
    core_instance1: bmg_72_324b883165919716
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp2: if ((core_name0 = "bmg_72_f580ae3be5511d30")) generate
    core_instance2: bmg_72_f580ae3be5511d30
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  comp3: if ((core_name0 = "bmg_72_3628803596b5ca22")) generate
    core_instance3: bmg_72_3628803596b5ca22
      port map (
        addra => core_addr,
        clka => clk,
        ena => core_ce,
        douta => core_data_out
                        );
  end generate;
  latency_test: if (latency > 1) generate
    reg: synth_reg
      generic map (
        width => c_width,
        latency => latency - 1
      )
      port map (
        i => core_data_out,
        ce => core_ce,
        clr => '0',
        clk => clk,
        o => data
      );
  end generate;
  latency_1: if (latency <= 1) generate
    data <= core_data_out;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_6e2bcf24f9 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_6e2bcf24f9;


architecture behavior of constant_6e2bcf24f9 is
begin
  op <= "10111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_54048c8b02 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54048c8b02;


architecture behavior of relational_54048c8b02 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xldpram_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    c_width_a: integer := 13;
    c_address_width_a: integer := 4;
    c_width_b: integer := 13;
    c_address_width_b: integer := 4;
    c_has_sinita: integer := 0;
    c_has_sinitb: integer := 0;
    latency: integer := 1
  );
  port (
    dina: in std_logic_vector(c_width_a - 1 downto 0);
    addra: in std_logic_vector(c_address_width_a - 1 downto 0);
    wea: in std_logic_vector(0 downto 0);
    a_ce: in std_logic;
    a_clk: in std_logic;
    rsta: in std_logic_vector(0 downto 0) := (others => '0');
    ena: in std_logic_vector(0 downto 0) := (others => '1');
    douta: out std_logic_vector(c_width_a - 1 downto 0);
    dinb: in std_logic_vector(c_width_b - 1 downto 0);
    addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
    web: in std_logic_vector(0 downto 0);
    b_ce: in std_logic;
    b_clk: in std_logic;
    rstb: in std_logic_vector(0 downto 0) := (others => '0');
    enb: in std_logic_vector(0 downto 0) := (others => '1');
    doutb: out std_logic_vector(c_width_b - 1 downto 0)
  );
end xldpram_wlan_phy_tx_pmd;
architecture behavior of xldpram_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer;
      latency: integer
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;

  signal core_addra: std_logic_vector(c_address_width_a - 1 downto 0);
  signal core_addrb: std_logic_vector(c_address_width_b - 1 downto 0);
  signal core_dina, core_douta, dly_douta:
    std_logic_vector(c_width_a - 1 downto 0);
  signal core_dinb, core_doutb, dly_doutb:
    std_logic_vector(c_width_b - 1 downto 0);
  signal core_wea, core_web: std_logic;
  signal core_a_ce, core_b_ce: std_logic;
  signal sinita, sinitb: std_logic;

  component bmg_72_7ec9033b751d2879
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_7ec9033b751d2879:
    component is true;
  attribute fpga_dont_touch of bmg_72_7ec9033b751d2879:
    component is "true";
  attribute box_type of bmg_72_7ec9033b751d2879:
    component  is "black_box";
  component bmg_72_da153342fc52049b
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_da153342fc52049b:
    component is true;
  attribute fpga_dont_touch of bmg_72_da153342fc52049b:
    component is "true";
  attribute box_type of bmg_72_da153342fc52049b:
    component  is "black_box";
  component bmg_72_41985f385eaacb3e
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_41985f385eaacb3e:
    component is true;
  attribute fpga_dont_touch of bmg_72_41985f385eaacb3e:
    component is "true";
  attribute box_type of bmg_72_41985f385eaacb3e:
    component  is "black_box";
  component bmg_72_376dc060ca4075f2
    port (
        addra: in std_logic_vector(c_address_width_a - 1 downto 0);
      addrb: in std_logic_vector(c_address_width_b - 1 downto 0);
      dina: in std_logic_vector(c_width_a - 1 downto 0);
      dinb: in std_logic_vector(c_width_b - 1 downto 0);
      clka: in std_logic;
      clkb: in std_logic;
      wea: in std_logic_vector(0 downto 0);
      web: in std_logic_vector(0 downto 0);
      ena: in std_logic;
      enb: in std_logic;
      douta: out std_logic_vector(c_width_a - 1 downto 0);
      doutb: out std_logic_vector(c_width_b - 1 downto 0)
     );
  end component;

  attribute syn_black_box of bmg_72_376dc060ca4075f2:
    component is true;
  attribute fpga_dont_touch of bmg_72_376dc060ca4075f2:
    component is "true";
  attribute box_type of bmg_72_376dc060ca4075f2:
    component  is "black_box";
begin
  core_addra <= addra;
  core_dina <= dina;
  douta <= dly_douta;
  core_wea <= wea(0);
  core_a_ce <= a_ce and ena(0);
  sinita <= rsta(0) and a_ce;

  core_addrb <= addrb;
  core_dinb <= dinb;
  doutb <= dly_doutb;
  core_web <= web(0);
  core_b_ce <= b_ce and enb(0);
  sinitb <= rstb(0) and b_ce;
  comp0: if ((core_name0 = "bmg_72_7ec9033b751d2879")) generate
    core_instance0: bmg_72_7ec9033b751d2879
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp1: if ((core_name0 = "bmg_72_da153342fc52049b")) generate
    core_instance1: bmg_72_da153342fc52049b
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp2: if ((core_name0 = "bmg_72_41985f385eaacb3e")) generate
    core_instance2: bmg_72_41985f385eaacb3e
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  comp3: if ((core_name0 = "bmg_72_376dc060ca4075f2")) generate
    core_instance3: bmg_72_376dc060ca4075f2
      port map (
          addra => core_addra,
        clka => a_clk,
        addrb => core_addrb,
        clkb => b_clk,
        dina => core_dina,
        wea(0) => core_wea,
        dinb => core_dinb,
        web(0) => core_web,
        ena => core_a_ce,
        enb => core_b_ce,
        douta => core_douta,
        doutb => core_doutb
      );
  end generate;
  latency_test: if (latency > 2) generate
    regA: synth_reg
      generic map (
        width => c_width_a,
        latency => latency - 2
      )
      port map (
        i => core_douta,
        ce => core_a_ce,
        clr => '0',
        clk => a_clk,
        o => dly_douta
      );
    regB: synth_reg
      generic map (
        width => c_width_b,
        latency => latency - 2
      )
      port map (
        i => core_doutb,
        ce => core_b_ce,
        clr => '0',
        clk => b_clk,
        o => dly_doutb
      );
  end generate;
  latency1: if (latency <= 2) generate
    dly_douta <= core_douta;
    dly_doutb <= core_doutb;
  end generate;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_1ece14600f is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((8 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_1ece14600f;


architecture behavior of concat_1ece14600f is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((8 - 1) downto 0);
  signal y_2_1_concat: unsigned((9 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_c6a9b6687e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_c6a9b6687e;


architecture behavior of concat_c6a9b6687e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((6 - 1) downto 0);
  signal y_2_1_concat: unsigned((7 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_4c449dd556 is
  port (
    op : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_4c449dd556;


architecture behavior of constant_4c449dd556 is
begin
  op <= "0000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8cac5f7cf5 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8cac5f7cf5;


architecture behavior of constant_8cac5f7cf5 is
begin
  op <= "011110010111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1bebc71bf9 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1bebc71bf9;


architecture behavior of constant_1bebc71bf9 is
begin
  op <= "100001101001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_92715f6857 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_92715f6857;


architecture behavior of constant_92715f6857 is
begin
  op <= "110101111000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9b9cbaee60 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9b9cbaee60;


architecture behavior of constant_9b9cbaee60 is
begin
  op <= "001010001000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_192c5da026 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    d3 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_192c5da026;


architecture behavior of mux_192c5da026 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal d3_1_33: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when "10" =>
        unregy_join_6_1 <= d2_1_30;
      when others =>
        unregy_join_6_1 <= d3_1_33;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8d143efc5e is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8d143efc5e;


architecture behavior of constant_8d143efc5e is
begin
  op <= "100011111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6c3ee657fa is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((9 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6c3ee657fa;


architecture behavior of relational_6c3ee657fa is
  signal a_1_31: unsigned((9 - 1) downto 0);
  signal b_1_34: unsigned((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_9779a5cf83 is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((10 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_9779a5cf83;


architecture behavior of concat_9779a5cf83 is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((9 - 1) downto 0);
  signal y_2_1_concat: unsigned((10 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_9127ce6619 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_9127ce6619;


architecture behavior of constant_9127ce6619 is
begin
  op <= "011111111111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_555e35158a is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_555e35158a;


architecture behavior of constant_555e35158a is
begin
  op <= "100111010100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_c0e78ca39c is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_c0e78ca39c;


architecture behavior of constant_c0e78ca39c is
begin
  op <= "110001001100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e3898a7c17 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e3898a7c17;


architecture behavior of constant_e3898a7c17 is
begin
  op <= "001110110100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_e054d850c5 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_e054d850c5;


architecture behavior of constant_e054d850c5 is
begin
  op <= "100000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_d3e8ce78bb is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_d3e8ce78bb;


architecture behavior of constant_d3e8ce78bb is
begin
  op <= "111011000100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_20bb1d9cec is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_20bb1d9cec;


architecture behavior of constant_20bb1d9cec is
begin
  op <= "000100111100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_044e9822dd is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_044e9822dd;


architecture behavior of constant_044e9822dd is
begin
  op <= "011000101100";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f3bb14635d is
  port (
    sel : in std_logic_vector((3 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    d3 : in std_logic_vector((12 - 1) downto 0);
    d4 : in std_logic_vector((12 - 1) downto 0);
    d5 : in std_logic_vector((12 - 1) downto 0);
    d6 : in std_logic_vector((12 - 1) downto 0);
    d7 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f3bb14635d;


architecture behavior of mux_f3bb14635d is
  signal sel_1_20: std_logic_vector((3 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal d3_1_33: std_logic_vector((12 - 1) downto 0);
  signal d4_1_36: std_logic_vector((12 - 1) downto 0);
  signal d5_1_39: std_logic_vector((12 - 1) downto 0);
  signal d6_1_42: std_logic_vector((12 - 1) downto 0);
  signal d7_1_45: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  d5_1_39 <= d5;
  d6_1_42 <= d6;
  d7_1_45 <= d7;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, d3_1_33, d4_1_36, d5_1_39, d6_1_42, d7_1_45, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "000" =>
        unregy_join_6_1 <= d0_1_24;
      when "001" =>
        unregy_join_6_1 <= d1_1_27;
      when "010" =>
        unregy_join_6_1 <= d2_1_30;
      when "011" =>
        unregy_join_6_1 <= d3_1_33;
      when "100" =>
        unregy_join_6_1 <= d4_1_36;
      when "101" =>
        unregy_join_6_1 <= d5_1_39;
      when "110" =>
        unregy_join_6_1 <= d6_1_42;
      when others =>
        unregy_join_6_1 <= d7_1_45;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_931d61fb72 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_931d61fb72;


architecture behavior of relational_931d61fb72 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_58c7454693 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_58c7454693;


architecture behavior of constant_58c7454693 is
begin
  op <= "100001100110";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_504d9a75aa is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_504d9a75aa;


architecture behavior of constant_504d9a75aa is
begin
  op <= "011110011010";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_fd28b32bf8 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_fd28b32bf8;


architecture behavior of constant_fd28b32bf8 is
begin
  op <= "000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_c3e1ddb86e is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_c3e1ddb86e;


architecture behavior of mux_c3e1ddb86e is
  signal sel_1_20: std_logic_vector((1 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_5c27e02321 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_5c27e02321;


architecture behavior of constant_5c27e02321 is
begin
  op <= "110000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4075671a27 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((6 - 1) downto 0);
    d1 : in std_logic_vector((9 - 1) downto 0);
    y : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4075671a27;


architecture behavior of mux_4075671a27 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((6 - 1) downto 0);
  signal d1_1_27: std_logic_vector((9 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((9 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= cast(d0_1_24, 0, 9, 0, xlUnsigned);
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_7b07120b87 is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7b07120b87;


architecture behavior of constant_7b07120b87 is
begin
  op <= "1000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_23065a6aa3 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_23065a6aa3;


architecture behavior of relational_23065a6aa3 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_14_3_rel <= a_1_31 /= b_1_34;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_1f05b15a2d is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_1f05b15a2d;


architecture behavior of constant_1f05b15a2d is
begin
  op <= "010101";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_330e503d71 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_330e503d71;


architecture behavior of constant_330e503d71 is
begin
  op <= "000111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_173d83e4a7 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_173d83e4a7;


architecture behavior of constant_173d83e4a7 is
begin
  op <= "111001";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_8207020ee3 is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8207020ee3;


architecture behavior of constant_8207020ee3 is
begin
  op <= "101011";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_e77c53f8bd is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_e77c53f8bd;


architecture behavior of logical_e77c53f8bd is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_4de2214a42 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_4de2214a42;


architecture behavior of mux_4de2214a42 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_47932db5b1 is
  port (
    a : in std_logic_vector((6 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_47932db5b1;


architecture behavior of relational_47932db5b1 is
  signal a_1_31: unsigned((6 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal result_16_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_16_3_rel <= a_1_31 < b_1_34;
  op <= boolean_to_vector(result_16_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_1834ac00b4 is
  port (
    a : in std_logic_vector((9 - 1) downto 0);
    b : in std_logic_vector((6 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_1834ac00b4;


architecture behavior of relational_1834ac00b4 is
  signal a_1_31: signed((9 - 1) downto 0);
  signal b_1_34: unsigned((6 - 1) downto 0);
  signal cast_12_17: signed((9 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_signed(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2s_cast(b_1_34, 0, 9, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity delay_0341f7be44 is
  port (
    d : in std_logic_vector((1 - 1) downto 0);
    q : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end delay_0341f7be44;


architecture behavior of delay_0341f7be44 is
  signal d_1_22: std_logic;
begin
  d_1_22 <= d(0);
  q <= std_logic_to_vector(d_1_22);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_011ca80190 is
  port (
    op : out std_logic_vector((7 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_011ca80190;


architecture behavior of constant_011ca80190 is
begin
  op <= "1011111";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_9a3978c602 is
  port (
    a : in std_logic_vector((7 - 1) downto 0);
    b : in std_logic_vector((7 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_9a3978c602;


architecture behavior of relational_9a3978c602 is
  signal a_1_31: unsigned((7 - 1) downto 0);
  signal b_1_34: unsigned((7 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_83e473517e is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((7 - 1) downto 0);
    y : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_83e473517e;


architecture behavior of concat_83e473517e is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((7 - 1) downto 0);
  signal y_2_1_concat: unsigned((8 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_2a9931b0e7 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_2a9931b0e7;


architecture behavior of constant_2a9931b0e7 is
begin
  op <= "101001011000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_40d4599892 is
  port (
    op : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_40d4599892;


architecture behavior of constant_40d4599892 is
begin
  op <= "010110101000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e6f5ee726b is
  port (
    in0 : in std_logic_vector((1 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e6f5ee726b;


architecture behavior of concat_e6f5ee726b is
  signal in0_1_23: unsigned((1 - 1) downto 0);
  signal in1_1_27: unsigned((1 - 1) downto 0);
  signal y_2_1_concat: unsigned((2 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= std_logic_vector_to_unsigned(in1);
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & unsigned_to_std_logic_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_33c9a0c803 is
  port (
    d0 : in std_logic_vector((2 - 1) downto 0);
    d1 : in std_logic_vector((2 - 1) downto 0);
    y : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_33c9a0c803;


architecture behavior of logical_33c9a0c803 is
  signal d0_1_24: std_logic_vector((2 - 1) downto 0);
  signal d1_1_27: std_logic_vector((2 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((2 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_e5a9964709 is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((12 - 1) downto 0);
    d1 : in std_logic_vector((12 - 1) downto 0);
    d2 : in std_logic_vector((12 - 1) downto 0);
    y : out std_logic_vector((12 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_e5a9964709;


architecture behavior of mux_e5a9964709 is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic_vector((12 - 1) downto 0);
  signal d1_1_27: std_logic_vector((12 - 1) downto 0);
  signal d2_1_30: std_logic_vector((12 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((12 - 1) downto 0);
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.conv_pkg.all;
entity xlfifogen_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    data_width: integer := -1;
    data_count_width: integer := -1;
    percent_full_width: integer := -1;
    has_ae : integer := 0;
    has_af : integer := 0
  );
  port (
    din: in std_logic_vector(data_width - 1 downto 0);
    we: in std_logic;
    we_ce: in std_logic;
    re: in std_logic;
    re_ce: in std_logic;
    rst: in std_logic;
    en: in std_logic;
    ce: in std_logic;
    clk: in std_logic;
    empty: out std_logic;
    full: out std_logic;
    percent_full: out std_logic_vector(percent_full_width - 1 downto 0);
    dcount: out std_logic_vector(data_count_width - 1 downto 0);
    ae: out std_logic;
    af: out std_logic;
    dout: out std_logic_vector(data_width - 1 downto 0)
  );
end xlfifogen_wlan_phy_tx_pmd ;
architecture behavior of xlfifogen_wlan_phy_tx_pmd is
  component fifo_fg92_6a1156e8dc43a711
    port (
      clk: in std_logic;
      srst: in std_logic;
      din: in std_logic_vector(data_width - 1 downto 0);
      wr_en: in std_logic;
      rd_en: in std_logic;
      dout: out std_logic_vector(data_width - 1 downto 0);
      full: out std_logic;
      empty: out std_logic;
      data_count: out std_logic_vector(data_count_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of fifo_fg92_6a1156e8dc43a711:
    component is true;
  attribute fpga_dont_touch of fifo_fg92_6a1156e8dc43a711:
    component is "true";
  attribute box_type of fifo_fg92_6a1156e8dc43a711:
    component  is "black_box";
  signal rd_en: std_logic;
  signal wr_en: std_logic;
  signal srst: std_logic;
  signal core_full: std_logic;
  signal core_dcount: std_logic_vector(data_count_width - 1 downto 0);
begin
  comp0: if ((core_name0 = "fifo_fg92_6a1156e8dc43a711")) generate
    core_instance0: fifo_fg92_6a1156e8dc43a711
      port map (
        clk => clk,
        srst => srst,
        din => din,
        wr_en => wr_en,
        rd_en => rd_en,
        dout => dout,
        full => core_full,
        empty => empty,
        data_count => core_dcount
      );
  end generate;

  modify_count: process(core_full, core_dcount) is
  begin
    if core_full = '1' then
      percent_full <= (others => '1');
    else
      percent_full <= core_dcount(data_count_width-1 downto data_count_width-percent_full_width);
    end if;
  end process modify_count;

  rd_en <= re and en and re_ce;
  wr_en <= we and en and we_ce;
  full <= core_full;
  srst <= rst and ce;
  dcount <= core_dcount;

  terminate_core_ae: if has_ae /= 1 generate
  begin
    ae <= '0';
  end generate terminate_core_ae;
  terminate_core_af: if has_af /= 1 generate
  begin
    af <= '0';
  end generate terminate_core_af;
end  behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_0512fd5e4c is
  port (
    op : out std_logic_vector((9 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0512fd5e4c;


architecture behavior of constant_0512fd5e4c is
begin
  op <= "100111111";
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.conv_pkg.all;
entity xlmult_wlan_phy_tx_pmd is
  generic (
    core_name0: string := "";
    a_width: integer := 4;
    a_bin_pt: integer := 2;
    a_arith: integer := xlSigned;
    b_width: integer := 4;
    b_bin_pt: integer := 1;
    b_arith: integer := xlSigned;
    p_width: integer := 8;
    p_bin_pt: integer := 2;
    p_arith: integer := xlSigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    extra_registers: integer := 0;
    c_a_width: integer := 7;
    c_b_width: integer := 7;
    c_type: integer := 0;
    c_a_type: integer := 0;
    c_b_type: integer := 0;
    c_pipelined: integer := 1;
    c_baat: integer := 4;
    multsign: integer := xlSigned;
    c_output_width: integer := 16
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    core_ce: in std_logic := '0';
    core_clr: in std_logic := '0';
    core_clk: in std_logic := '0';
    rst: in std_logic_vector(rst_width - 1 downto 0);
    en: in std_logic_vector(en_width - 1 downto 0);
    p: out std_logic_vector(p_width - 1 downto 0)
  );
end xlmult_wlan_phy_tx_pmd;
architecture behavior of xlmult_wlan_phy_tx_pmd is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component mult_11_2_f2bb5a57782af7d9
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of mult_11_2_f2bb5a57782af7d9:
    component is true;
  attribute fpga_dont_touch of mult_11_2_f2bb5a57782af7d9:
    component is "true";
  attribute box_type of mult_11_2_f2bb5a57782af7d9:
    component  is "black_box";
  component mult_11_2_414c0fa5acc33f35
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;

  attribute syn_black_box of mult_11_2_414c0fa5acc33f35:
    component is true;
  attribute fpga_dont_touch of mult_11_2_414c0fa5acc33f35:
    component is "true";
  attribute box_type of mult_11_2_414c0fa5acc33f35:
    component  is "black_box";
  signal tmp_a: std_logic_vector(c_a_width - 1 downto 0);
  signal conv_a: std_logic_vector(c_a_width - 1 downto 0);
  signal tmp_b: std_logic_vector(c_b_width - 1 downto 0);
  signal conv_b: std_logic_vector(c_b_width - 1 downto 0);
  signal tmp_p: std_logic_vector(c_output_width - 1 downto 0);
  signal conv_p: std_logic_vector(p_width - 1 downto 0);
  -- synopsys translate_off
  signal real_a, real_b, real_p: real;
  -- synopsys translate_on
  signal rfd: std_logic;
  signal rdy: std_logic;
  signal nd: std_logic;
  signal internal_ce: std_logic;
  signal internal_clr: std_logic;
  signal internal_core_ce: std_logic;
begin
-- synopsys translate_off
-- synopsys translate_on
  internal_ce <= ce and en(0);
  internal_core_ce <= core_ce and en(0);
  internal_clr <= (clr or rst(0)) and ce;
  nd <= internal_ce;
  input_process:  process (a,b)
  begin
    tmp_a <= zero_ext(a, c_a_width);
    tmp_b <= zero_ext(b, c_b_width);
  end process;
  output_process: process (tmp_p)
  begin
    conv_p <= convert_type(tmp_p, c_output_width, a_bin_pt+b_bin_pt, multsign,
                           p_width, p_bin_pt, p_arith, quantization, overflow);
  end process;
  comp0: if ((core_name0 = "mult_11_2_f2bb5a57782af7d9")) generate
    core_instance0: mult_11_2_f2bb5a57782af7d9
      port map (
        a => tmp_a,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  comp1: if ((core_name0 = "mult_11_2_414c0fa5acc33f35")) generate
    core_instance1: mult_11_2_414c0fa5acc33f35
      port map (
        a => tmp_a,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  latency_gt_0: if (extra_registers > 0) generate
    reg: synth_reg
      generic map (
        width => p_width,
        latency => extra_registers
      )
      port map (
        i => conv_p,
        ce => internal_ce,
        clr => internal_clr,
        clk => clk,
        o => p
      );
  end generate;
  latency_eq_0: if (extra_registers = 0) generate
    p <= conv_p;
  end generate;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_a54904b290 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((16 - 1) downto 0);
    d1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_a54904b290;


architecture behavior of mux_a54904b290 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((16 - 1) downto 0);
  signal d1_1_27: std_logic_vector((16 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((16 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_bfe1d4f686 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((16 - 1) downto 0);
    d1 : in std_logic_vector((16 - 1) downto 0);
    y : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_bfe1d4f686;


architecture behavior of mux_bfe1d4f686 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((16 - 1) downto 0);
  signal d1_1_27: std_logic_vector((16 - 1) downto 0);
  type array_type_pipe_16_22 is array (0 to (1 - 1)) of std_logic_vector((16 - 1) downto 0);
  signal pipe_16_22: array_type_pipe_16_22 := (
    0 => "0000000000000000");
  signal pipe_16_22_front_din: std_logic_vector((16 - 1) downto 0);
  signal pipe_16_22_back: std_logic_vector((16 - 1) downto 0);
  signal pipe_16_22_push_front_pop_back_en: std_logic;
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((16 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  pipe_16_22_back <= pipe_16_22(0);
  proc_pipe_16_22: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (pipe_16_22_push_front_pop_back_en = '1')) then
        pipe_16_22(0) <= pipe_16_22_front_din;
      end if;
    end if;
  end process proc_pipe_16_22;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  pipe_16_22_front_din <= unregy_join_6_1;
  pipe_16_22_push_front_pop_back_en <= '1';
  y <= pipe_16_22_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_6dad3a03fc is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_6dad3a03fc;


architecture behavior of relational_6dad3a03fc is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_12_17: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 8, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity concat_e25f797841 is
  port (
    in0 : in std_logic_vector((31 - 1) downto 0);
    in1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end concat_e25f797841;


architecture behavior of concat_e25f797841 is
  signal in0_1_23: unsigned((31 - 1) downto 0);
  signal in1_1_27: boolean;
  signal y_2_1_concat: unsigned((32 - 1) downto 0);
begin
  in0_1_23 <= std_logic_vector_to_unsigned(in0);
  in1_1_27 <= ((in1) = "1");
  y_2_1_concat <= std_logic_vector_to_unsigned(unsigned_to_std_logic_vector(in0_1_23) & boolean_to_vector(in1_1_27));
  y <= unsigned_to_std_logic_vector(y_2_1_concat);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_bc7a810978 is
  port (
    op : out std_logic_vector((31 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_bc7a810978;


architecture behavior of constant_bc7a810978 is
begin
  op <= "0000000000000000000000000000000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity reinterpret_ddc3ebdd7c is
  port (
    input_port : in std_logic_vector((16 - 1) downto 0);
    output_port : out std_logic_vector((16 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end reinterpret_ddc3ebdd7c;


architecture behavior of reinterpret_ddc3ebdd7c is
  signal input_port_1_40: unsigned((16 - 1) downto 0);
begin
  input_port_1_40 <= std_logic_vector_to_unsigned(input_port);
  output_port <= unsigned_to_std_logic_vector(input_port_1_40);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_899cf9b568 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    d3 : in std_logic_vector((1 - 1) downto 0);
    d4 : in std_logic_vector((1 - 1) downto 0);
    en : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_899cf9b568;


architecture behavior of logical_899cf9b568 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal d3_1_33: std_logic_vector((1 - 1) downto 0);
  signal d4_1_36: std_logic_vector((1 - 1) downto 0);
  signal en_1_39: std_logic;
  type array_type_latency_pipe_5_26 is array (0 to (1 - 1)) of std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26: array_type_latency_pipe_5_26 := (
    0 => "0");
  signal latency_pipe_5_26_front_din: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_back: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_5_26_push_front_pop_back_en: std_logic;
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_shift_join_7_1: std_logic_vector((1 - 1) downto 0);
  signal latency_pipe_shift_join_7_1_en: std_logic;
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  d3_1_33 <= d3;
  d4_1_36 <= d4;
  en_1_39 <= en(0);
  latency_pipe_5_26_back <= latency_pipe_5_26(0);
  proc_latency_pipe_5_26: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (latency_pipe_5_26_push_front_pop_back_en = '1')) then
        latency_pipe_5_26(0) <= latency_pipe_5_26_front_din;
      end if;
    end if;
  end process proc_latency_pipe_5_26;
  fully_2_1_bit <= d0_1_24 xor d1_1_27 xor d2_1_30 xor d3_1_33 xor d4_1_36;
  proc_if_7_1: process (en_1_39, fully_2_1_bit)
  is
  begin
    if en_1_39 = '1' then
      latency_pipe_shift_join_7_1_en <= '1';
    else 
      latency_pipe_shift_join_7_1_en <= '0';
    end if;
    latency_pipe_shift_join_7_1 <= fully_2_1_bit;
  end process proc_if_7_1;
  latency_pipe_5_26_front_din <= latency_pipe_shift_join_7_1;
  latency_pipe_5_26_push_front_pop_back_en <= latency_pipe_shift_join_7_1_en;
  y <= latency_pipe_5_26_back;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity constant_3a9a3daeb9 is
  port (
    op : out std_logic_vector((2 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_3a9a3daeb9;


architecture behavior of constant_3a9a3daeb9 is
begin
  op <= "11";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_5f1eb17108 is
  port (
    a : in std_logic_vector((2 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_5f1eb17108;


architecture behavior of relational_5f1eb17108 is
  signal a_1_31: unsigned((2 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_706b9eb7ce is
  port (
    a : in std_logic_vector((3 - 1) downto 0);
    b : in std_logic_vector((2 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_706b9eb7ce;


architecture behavior of relational_706b9eb7ce is
  signal a_1_31: unsigned((3 - 1) downto 0);
  signal b_1_34: unsigned((2 - 1) downto 0);
  signal cast_12_17: unsigned((3 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 3, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_472286caed is
  port (
    sel : in std_logic_vector((2 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_472286caed;


architecture behavior of mux_472286caed is
  signal sel_1_20: std_logic_vector((2 - 1) downto 0);
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal d2_1_30: std_logic;
  signal unregy_join_6_1: std_logic;
begin
  sel_1_20 <= sel;
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  d2_1_30 <= d2(0);
  proc_switch_6_1: process (d0_1_24, d1_1_27, d2_1_30, sel_1_20)
  is
  begin
    case sel_1_20 is 
      when "00" =>
        unregy_join_6_1 <= d0_1_24;
      when "01" =>
        unregy_join_6_1 <= d1_1_27;
      when others =>
        unregy_join_6_1 <= d2_1_30;
    end case;
  end process proc_switch_6_1;
  y <= std_logic_to_vector(unregy_join_6_1);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_9d76333483 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_9d76333483;


architecture behavior of logical_9d76333483 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 xor d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_7b6bf7e572 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    d2 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_7b6bf7e572;


architecture behavior of logical_7b6bf7e572 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal d2_1_30: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  fully_2_1_bit <= d0_1_24 and d1_1_27 and d2_1_30;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_112ed141f4 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_112ed141f4;


architecture behavior of mux_112ed141f4 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((1 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity relational_7bfd319389 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_7bfd319389;


architecture behavior of relational_7bfd319389 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_18_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_18_3_rel <= a_1_31 > b_1_34;
  op <= boolean_to_vector(result_18_3_rel);
end behavior;


-------------------------------------------------------------------
-- System Generator version 14.3 VHDL source file.
--
-- Copyright(C) 2012 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2012 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
entity xlusamp is
    generic (
             d_width      : integer := 5;
             d_bin_pt     : integer := 2;
             d_arith      : integer := xlUnsigned;
             q_width      : integer := 5;
             q_bin_pt     : integer := 2;
             q_arith      : integer := xlUnsigned;
             en_width     : integer := 1;
             en_bin_pt    : integer := 0;
             en_arith     : integer := xlUnsigned;
             sampling_ratio     : integer := 2;
             latency      : integer := 1;
             copy_samples : integer := 0);
    port (
          d        : in std_logic_vector (d_width-1 downto 0);
          src_clk  : in std_logic;
          src_ce   : in std_logic;
          src_clr  : in std_logic;
          dest_clk : in std_logic;
          dest_ce  : in std_logic;
          dest_clr : in std_logic;
          en       : in std_logic_vector(en_width-1 downto 0);
          q        : out std_logic_vector (q_width-1 downto 0)
         );
end xlusamp;
architecture struct of xlusamp is
    component synth_reg
      generic (
        width: integer := 16;
        latency: integer := 5
      );
      port (
        i: in std_logic_vector(width - 1 downto 0);
        ce: in std_logic;
        clr: in std_logic;
        clk: in std_logic;
        o: out std_logic_vector(width - 1 downto 0)
      );
    end component;
    component FDSE
        port (q  : out   std_ulogic;
              d  : in    std_ulogic;
              c  : in    std_ulogic;
              s  : in    std_ulogic;
              ce : in    std_ulogic);
    end component;
    attribute syn_black_box of FDSE : component is true;
    attribute fpga_dont_touch of FDSE : component is "true";
    signal zero    : std_logic_vector (d_width-1 downto 0);
    signal mux_sel : std_logic;
    signal sampled_d  : std_logic_vector (d_width-1 downto 0);
    signal internal_ce : std_logic;
begin
   sel_gen : FDSE
                port map (q  => mux_sel,
                        d  => src_ce,
            c  => src_clk,
            s  => src_clr,
            ce => dest_ce);
  internal_ce <= src_ce and en(0);
  copy_samples_false : if (copy_samples = 0) generate
      zero <= (others => '0');
      gen_q_cp_smpls_0_and_lat_0: if (latency = 0) generate
        cp_smpls_0_and_lat_0: process (mux_sel, d, zero)
        begin
          if (mux_sel = '1') then
            q <= d;
          else
            q <= zero;
          end if;
        end process cp_smpls_0_and_lat_0;
      end generate;
      gen_q_cp_smpls_0_and_lat_gt_0: if (latency > 0) generate
        sampled_d_reg: synth_reg
          generic map (
            width => d_width,
            latency => latency
          )
          port map (
            i => d,
            ce => internal_ce,
            clr => src_clr,
            clk => src_clk,
            o => sampled_d
          );

        gen_q_check_mux_sel: process (mux_sel, sampled_d, zero)
        begin
          if (mux_sel = '1') then
            q <= sampled_d;
          else
            q <= zero;
          end if;
        end process gen_q_check_mux_sel;
      end generate;
   end generate;
   copy_samples_true : if (copy_samples = 1) generate
     gen_q_cp_smpls_1_and_lat_0: if (latency = 0) generate
       q <= d;
     end generate;
     gen_q_cp_smpls_1_and_lat_gt_0: if (latency > 0) generate
       q <= sampled_d;
       sampled_d_reg2: synth_reg
         generic map (
           width => d_width,
           latency => latency
         )
         port map (
           i => d,
           ce => internal_ce,
           clr => src_clr,
           clk => src_clk,
           o => sampled_d
         );
     end generate;
   end generate;
end architecture struct;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity mux_f9c0f11a18 is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((4 - 1) downto 0);
    d1 : in std_logic_vector((4 - 1) downto 0);
    y : out std_logic_vector((4 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_f9c0f11a18;


architecture behavior of mux_f9c0f11a18 is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((4 - 1) downto 0);
  signal d1_1_27: std_logic_vector((4 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((4 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.conv_pkg.all;

entity logical_938d99ac11 is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_938d99ac11;


architecture behavior of logical_938d99ac11 is
  signal d0_1_24: std_logic_vector((1 - 1) downto 0);
  signal d1_1_27: std_logic_vector((1 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((1 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  fully_2_1_bit <= d0_1_24 and d1_1_27;
  y <= fully_2_1_bit;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Addr Gen"

entity addr_gen_entity_b968174b41 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    signal_length: in std_logic_vector(11 downto 0); 
    tx_reset: in std_logic; 
    bit_mem_addr: out std_logic_vector(14 downto 0); 
    data: out std_logic; 
    fcs: out std_logic; 
    pad: out std_logic; 
    ppdu_tail_done: out std_logic; 
    signal_x0: out std_logic; 
    tail: out std_logic
  );
end addr_gen_entity_b968174b41;

architecture structural of addr_gen_entity_b968174b41 is
  signal accumulator_q_net_x0: std_logic_vector(14 downto 0);
  signal addsub1_s_net: std_logic_vector(11 downto 0);
  signal addsub_s_net: std_logic_vector(11 downto 0);
  signal assert_dout_net: std_logic_vector(14 downto 0);
  signal b_16_5_y_net: std_logic_vector(11 downto 0);
  signal byte_addr_y_net: std_logic_vector(11 downto 0);
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(3 downto 0);
  signal constant3_op_net: std_logic_vector(4 downto 0);
  signal constant4_op_net: std_logic_vector(4 downto 0);
  signal constant5_op_net: std_logic_vector(5 downto 0);
  signal constant6_op_net: std_logic_vector(3 downto 0);
  signal constant7_op_net: std_logic_vector(4 downto 0);
  signal constant8_op_net: std_logic_vector(2 downto 0);
  signal constant9_op_net: std_logic_vector(2 downto 0);
  signal convert1_dout_net: std_logic;
  signal convert_dout_net: std_logic;
  signal delay3_q_net_x0: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal inverter4_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical4_y_net: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net_x0: std_logic;
  signal mux_y_net: std_logic_vector(4 downto 0);
  signal register_q_net_x0: std_logic;
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal relational3_op_net: std_logic;
  signal relational4_op_net: std_logic;
  signal relational5_op_net: std_logic;
  signal relational6_op_net_x0: std_logic;
  signal relational_op_net: std_logic;
  signal tail_bit_count_op_net: std_logic_vector(2 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  register_q_net_x0 <= en;
  b_16_5_y_net <= signal_length;
  logical_y_net_x0 <= tx_reset;
  bit_mem_addr <= accumulator_q_net_x0;
  data <= logical2_y_net_x0;
  fcs <= logical1_y_net_x0;
  pad <= relational6_op_net_x0;
  ppdu_tail_done <= delay3_q_net_x0;
  signal_x0 <= logical5_y_net_x0;
  tail <= logical3_y_net_x0;

  accumulator: entity work.accum_a764547d38
    port map (
      b => mux_y_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q => accumulator_q_net_x0
    );

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 12,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 4,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 13,
      core_name0 => "addsb_11_0_913f4bce6842c815",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 13,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 12
    )
    port map (
      a => byte_addr_y_net,
      b => constant6_op_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  addsub1: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 12,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 3,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 13,
      core_name0 => "addsb_11_0_913f4bce6842c815",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 13,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 12
    )
    port map (
      a => b_16_5_y_net,
      b => constant8_op_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => addsub1_s_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 15,
      dout_width => 15
    )
    port map (
      din => accumulator_q_net_x0,
      dout => assert_dout_net
    );

  byte_addr: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 14,
      x_width => 15,
      y_width => 12
    )
    port map (
      x => accumulator_q_net_x0,
      y => byte_addr_y_net
    );

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => relational_op_net,
      in1(0) => relational1_op_net,
      y => concat_y_net
    );

  constant1: entity work.constant_a7e2bb9e12
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_a629aefb53
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_f5633478bf
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_07db25d611
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_ef95fb0eb4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_145086465d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  constant7: entity work.constant_bc74ae1a6c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net
    );

  constant8: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net
    );

  constant9: entity work.constant_4e64dfaf34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant9_op_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => logical_y_net_x0,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => register_q_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => relational6_op_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x0
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip(0) => relational2_op_net,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip(0) => relational4_op_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip(0) => relational6_op_net_x0,
      op(0) => inverter3_op_net
    );

  inverter4: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip(0) => relational6_op_net_x0,
      op(0) => inverter4_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter2_op_net,
      d1(0) => relational3_op_net,
      y(0) => logical1_y_net_x0
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational4_op_net,
      d1(0) => inverter1_op_net,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational5_op_net,
      d1(0) => inverter3_op_net,
      y(0) => logical3_y_net_x0
    );

  logical4: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational5_op_net,
      d1(0) => convert1_dout_net,
      d2(0) => inverter4_op_net,
      y(0) => logical4_y_net
    );

  logical5: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => relational2_op_net,
      y(0) => logical5_y_net_x0
    );

  mux: entity work.mux_4a20039e59
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant1_op_net,
      d1 => constant2_op_net,
      d2 => constant3_op_net,
      sel => concat_y_net,
      y => mux_y_net
    );

  relational: entity work.relational_ec1b27521c
    port map (
      a => assert_dout_net,
      b => constant5_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity work.relational_37ecee0ab7
    port map (
      a => assert_dout_net,
      b => constant4_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_eed86727d9
    port map (
      a => accumulator_q_net_x0,
      b => constant7_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  relational3: entity work.relational_70fbe7d900
    port map (
      a => addsub_s_net,
      b => b_16_5_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  relational4: entity work.relational_70fbe7d900
    port map (
      a => addsub_s_net,
      b => addsub1_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  relational5: entity work.relational_b307c14bb5
    port map (
      a => addsub_s_net,
      b => b_16_5_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net
    );

  relational6: entity work.relational_07bde14ec5
    port map (
      a => tail_bit_count_op_net,
      b => constant9_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational6_op_net_x0
    );

  tail_bit_count: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 6,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_bcc28bfecf25caff",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 3
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => logical4_y_net,
      rst(0) => logical_y_net_x0,
      op => tail_bit_count_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/BRAM IF 64b"

entity bram_if_64b_entity_672a3af05d is
  port (
    bit_addr: in std_logic_vector(14 downto 0); 
    bram_din: in std_logic_vector(63 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    regtx_pkt_buf_addr_offset: in std_logic_vector(7 downto 0); 
    tx_pkt_buf_sel: in std_logic_vector(3 downto 0); 
    concat_x0: out std_logic_vector(31 downto 0); 
    constant1_x0: out std_logic; 
    constant2_x0: out std_logic; 
    constant7_x0: out std_logic_vector(63 downto 0); 
    constant8_x0: out std_logic_vector(7 downto 0); 
    x64b_data: out std_logic_vector(63 downto 0)
  );
end bram_if_64b_entity_672a3af05d;

architecture structural of bram_if_64b_entity_672a3af05d is
  signal accumulator_q_net_x1: std_logic_vector(14 downto 0);
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal b_23_16_y_net_x0: std_logic_vector(7 downto 0);
  signal bram_din_net_x0: std_logic_vector(63 downto 0);
  signal ce_1_sg_x1: std_logic;
  signal clk_1_sg_x1: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant1_op_net_x0: std_logic;
  signal constant2_op_net_x0: std_logic;
  signal constant3_op_net: std_logic_vector(2 downto 0);
  signal constant4_op_net: std_logic_vector(15 downto 0);
  signal constant7_op_net_x0: std_logic_vector(63 downto 0);
  signal constant8_op_net_x0: std_logic_vector(7 downto 0);
  signal mux_y_net_x0: std_logic_vector(3 downto 0);
  signal simulation_multiplexer_dout_net_x0: std_logic_vector(63 downto 0);
  signal x9msb_y_net: std_logic_vector(8 downto 0);

begin
  accumulator_q_net_x1 <= bit_addr;
  bram_din_net_x0 <= bram_din;
  ce_1_sg_x1 <= ce_1;
  clk_1_sg_x1 <= clk_1;
  b_23_16_y_net_x0 <= regtx_pkt_buf_addr_offset;
  mux_y_net_x0 <= tx_pkt_buf_sel;
  concat_x0 <= concat_y_net_x0;
  constant1_x0 <= constant1_op_net_x0;
  constant2_x0 <= constant2_op_net_x0;
  constant7_x0 <= constant7_op_net_x0;
  constant8_x0 <= constant8_op_net_x0;
  x64b_data <= simulation_multiplexer_dout_net_x0;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 9,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 8,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 10,
      core_name0 => "addsb_11_0_73986f767e994888",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 10,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => x9msb_y_net,
      b => b_23_16_y_net_x0,
      ce => ce_1_sg_x1,
      clk => clk_1_sg_x1,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  concat: entity work.concat_c5804edea5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant4_op_net,
      in1 => mux_y_net_x0,
      in2 => addsub_s_net,
      in3 => constant3_op_net,
      y => concat_y_net_x0
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net_x0
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net_x0
    );

  constant3: entity work.constant_822933f89b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_9f5572ba51
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant7: entity work.constant_c4c603edf2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net_x0
    );

  constant8: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net_x0
    );

  simulation_multiplexer: entity work.xlpassthrough
    generic map (
      din_width => 64,
      dout_width => 64
    )
    port map (
      din => bram_din_net_x0,
      dout => simulation_multiplexer_dout_net_x0
    );

  x9msb: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 14,
      x_width => 15,
      y_width => 9
    )
    port map (
      x => accumulator_q_net_x1,
      y => x9msb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Bit Per Sym Counter/Osc"

entity osc_entity_d1c47b8b4b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    q: out std_logic
  );
end osc_entity_d1c47b8b4b;

architecture structural of osc_entity_d1c47b8b4b is
  signal assert_dout_net: std_logic;
  signal ce_1_sg_x2: std_logic;
  signal clk_1_sg_x2: std_logic;
  signal inverter1_op_net: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register_q_net_x1: std_logic;

begin
  ce_1_sg_x2 <= ce_1;
  clk_1_sg_x2 <= clk_1;
  register2_q_net_x0 <= en;
  logical3_y_net_x0 <= rst;
  q <= register_q_net_x1;

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register_q_net_x1,
      dout(0) => assert_dout_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x2,
      clk => clk_1_sg_x2,
      clr => '0',
      ip(0) => assert_dout_net,
      op(0) => inverter1_op_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x2,
      clk => clk_1_sg_x2,
      d(0) => inverter1_op_net,
      en(0) => register2_q_net_x0,
      rst(0) => logical3_y_net_x0,
      q(0) => register_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Bit Per Sym Counter/Posedge1"

entity posedge1_entity_9966c21e4f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end posedge1_entity_9966c21e4f;

architecture structural of posedge1_entity_9966c21e4f is
  signal ce_1_sg_x3: std_logic;
  signal clk_1_sg_x3: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;

begin
  ce_1_sg_x3 <= ce_1;
  clk_1_sg_x3 <= clk_1;
  logical1_y_net_x1 <= d;
  q <= logical1_y_net_x2;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      d(0) => logical1_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x3,
      clk => clk_1_sg_x3,
      clr => '0',
      ip(0) => delay_q_net,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Bit Per Sym Counter/S-R Latch1"

entity s_r_latch1_entity_7106e36b8f is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    r: in std_logic; 
    s: in std_logic; 
    q: out std_logic
  );
end s_r_latch1_entity_7106e36b8f;

architecture structural of s_r_latch1_entity_7106e36b8f is
  signal ce_1_sg_x4: std_logic;
  signal clk_1_sg_x4: std_logic;
  signal constant1_op_net: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;

begin
  ce_1_sg_x4 <= ce_1;
  clk_1_sg_x4 <= clk_1;
  logical2_y_net_x0 <= r;
  logical1_y_net_x3 <= s;
  q <= register2_q_net_x1;

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      din(0) => logical2_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      clr => '0',
      din(0) => logical1_y_net_x3,
      en => "1",
      dout(0) => convert2_dout_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x4,
      clk => clk_1_sg_x4,
      d(0) => constant1_op_net,
      en(0) => convert2_dout_net,
      rst(0) => convert1_dout_net,
      q(0) => register2_q_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Bit Per Sym Counter"

entity bit_per_sym_counter_entity_be13008040 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_n_dbps: in std_logic_vector(8 downto 0); 
    start_sym: in std_logic; 
    tx_reset: in std_logic; 
    last_bit_in_sym: out std_logic; 
    load_bit: out std_logic
  );
end bit_per_sym_counter_entity_be13008040;

architecture structural of bit_per_sym_counter_entity_be13008040 is
  signal ce_1_sg_x6: std_logic;
  signal clk_1_sg_x6: std_logic;
  signal constant2_op_net: std_logic_vector(4 downto 0);
  signal convert3_dout_net_x0: std_logic_vector(8 downto 0);
  signal inverter_op_net_x1: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical_y_net_x2: std_logic;
  signal mux_y_net: std_logic_vector(8 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register_q_net_x2: std_logic;
  signal relational2_op_net: std_logic;
  signal sym_data_bit_count_op_net: std_logic_vector(8 downto 0);

begin
  ce_1_sg_x6 <= ce_1;
  clk_1_sg_x6 <= clk_1;
  convert3_dout_net_x0 <= data_n_dbps;
  logical1_y_net_x2 <= start_sym;
  logical_y_net_x2 <= tx_reset;
  last_bit_in_sym <= inverter_op_net_x1;
  load_bit <= register_q_net_x2;

  constant2: entity work.constant_bc74ae1a6c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      ip(0) => relational2_op_net,
      op(0) => inverter_op_net_x1
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net_x1,
      d1(0) => logical_y_net_x2,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x2,
      d1(0) => inverter_op_net_x1,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x2,
      d1(0) => inverter_op_net_x1,
      y(0) => logical3_y_net_x0
    );

  mux: entity work.mux_129040d58e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => convert3_dout_net_x0,
      sel(0) => register2_q_net_x0,
      y => mux_y_net
    );

  osc_d1c47b8b4b: entity work.osc_entity_d1c47b8b4b
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      en => register2_q_net_x1,
      rst => logical3_y_net_x0,
      q => register_q_net_x2
    );

  posedge1_9966c21e4f: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      d => logical1_y_net_x2,
      q => logical1_y_net_x3
    );

  relational2: entity work.relational_82fb466a8b
    port map (
      a => sym_data_bit_count_op_net,
      b => mux_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  s_r_latch1_7106e36b8f: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      r => logical2_y_net_x0,
      s => logical1_y_net_x3,
      q => register2_q_net_x1
    );

  s_r_latch2_b16421a885: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x6,
      clk_1 => clk_1_sg_x6,
      r => logical_y_net_x2,
      s => inverter_op_net_x1,
      q => register2_q_net_x0
    );

  sym_data_bit_count: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_36e2bb554c95560d",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x6,
      clk => clk_1_sg_x6,
      clr => '0',
      en(0) => register_q_net_x2,
      rst(0) => logical1_y_net,
      op => sym_data_bit_count_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/Bit Sel"

entity bit_sel_entity_2c3a4baaeb is
  port (
    b: in std_logic_vector(7 downto 0); 
    b_sel: in std_logic_vector(2 downto 0); 
    b_x0: out std_logic
  );
end bit_sel_entity_2c3a4baaeb;

architecture structural of bit_sel_entity_2c3a4baaeb is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b4_y_net: std_logic;
  signal b5_y_net: std_logic;
  signal b6_y_net: std_logic;
  signal b7_y_net: std_logic;
  signal mux_y_net_x1: std_logic_vector(7 downto 0);
  signal mux_y_net_x2: std_logic;
  signal x3lsb_y_net_x0: std_logic_vector(2 downto 0);

begin
  mux_y_net_x1 <= b;
  x3lsb_y_net_x0 <= b_sel;
  b_x0 <= mux_y_net_x2;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x1,
      y(0) => b7_y_net
    );

  mux: entity work.mux_b0082e75ff
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => b0_y_net,
      d1(0) => b1_y_net,
      d2(0) => b2_y_net,
      d3(0) => b3_y_net,
      d4(0) => b4_y_net,
      d5(0) => b5_y_net,
      d6(0) => b6_y_net,
      d7(0) => b7_y_net,
      sel => x3lsb_y_net_x0,
      y(0) => mux_y_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/Byte Sel"

entity byte_sel_entity_1b5e475260 is
  port (
    b_sel: in std_logic_vector(2 downto 0); 
    x64b: in std_logic_vector(63 downto 0); 
    b: out std_logic_vector(7 downto 0)
  );
end byte_sel_entity_1b5e475260;

architecture structural of byte_sel_entity_1b5e475260 is
  signal b0_y_net: std_logic_vector(7 downto 0);
  signal b1_y_net: std_logic_vector(7 downto 0);
  signal b2_y_net: std_logic_vector(7 downto 0);
  signal b3_y_net: std_logic_vector(7 downto 0);
  signal b4_y_net: std_logic_vector(7 downto 0);
  signal b5_y_net: std_logic_vector(7 downto 0);
  signal b6_y_net: std_logic_vector(7 downto 0);
  signal b7_y_net: std_logic_vector(7 downto 0);
  signal mux_y_net_x2: std_logic_vector(2 downto 0);
  signal mux_y_net_x3: std_logic_vector(63 downto 0);
  signal mux_y_net_x4: std_logic_vector(7 downto 0);

begin
  mux_y_net_x2 <= b_sel;
  mux_y_net_x3 <= x64b;
  b <= mux_y_net_x4;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 32,
      new_msb => 39,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 40,
      new_msb => 47,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 48,
      new_msb => 55,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 56,
      new_msb => 63,
      x_width => 64,
      y_width => 8
    )
    port map (
      x => mux_y_net_x3,
      y => b7_y_net
    );

  mux: entity work.mux_c762ea476a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b0_y_net,
      d1 => b1_y_net,
      d2 => b2_y_net,
      d3 => b3_y_net,
      d4 => b4_y_net,
      d5 => b5_y_net,
      d6 => b6_y_net,
      d7 => b7_y_net,
      sel => mux_y_net_x2,
      y => mux_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/Byte sel"

entity byte_sel_entity_3a45df7438 is
  port (
    bit_ind: in std_logic_vector(14 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    src_sel: in std_logic_vector(1 downto 0); 
    tx_reset: in std_logic; 
    sel: out std_logic_vector(2 downto 0)
  );
end byte_sel_entity_3a45df7438;

architecture structural of byte_sel_entity_3a45df7438 is
  signal ce_1_sg_x8: std_logic;
  signal clk_1_sg_x8: std_logic;
  signal concat_y_net_x0: std_logic_vector(1 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(2 downto 0);
  signal counter_op_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x0: std_logic_vector(14 downto 0);
  signal delay_q_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical_y_net_x3: std_logic;
  signal lsb_y_net: std_logic;
  signal mux_y_net_x3: std_logic_vector(2 downto 0);
  signal relational3_op_net: std_logic;
  signal x3lsb_3_y_net: std_logic_vector(2 downto 0);
  signal x3lsb_y_net: std_logic_vector(2 downto 0);

begin
  delay1_q_net_x0 <= bit_ind;
  ce_1_sg_x8 <= ce_1;
  clk_1_sg_x8 <= clk_1;
  concat_y_net_x0 <= src_sel;
  logical_y_net_x3 <= tx_reset;
  sel <= mux_y_net_x3;

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_1d6ad1c713
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_6454489cfe866515",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x8,
      clk => clk_1_sg_x8,
      clr => '0',
      en(0) => logical1_y_net_x2,
      rst(0) => logical_y_net_x3,
      op => counter_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x8,
      clk => clk_1_sg_x8,
      d(0) => relational3_op_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  logical1: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => lsb_y_net,
      d1(0) => relational3_op_net,
      d2(0) => delay_q_net,
      y(0) => logical1_y_net_x1
    );

  lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => concat_y_net_x0,
      y(0) => lsb_y_net
    );

  mux: entity work.mux_a10351e9f3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => x3lsb_3_y_net,
      d1 => counter_op_net,
      d2 => constant1_op_net,
      sel => concat_y_net_x0,
      y => mux_y_net_x3
    );

  posedge_5f4bf4b001: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x8,
      clk_1 => clk_1_sg_x8,
      d => logical1_y_net_x1,
      q => logical1_y_net_x2
    );

  relational3: entity work.relational_8fc7f5539b
    port map (
      a => x3lsb_y_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  x3lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 15,
      y_width => 3
    )
    port map (
      x => delay1_q_net_x0,
      y => x3lsb_y_net
    );

  x3lsb_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 5,
      x_width => 15,
      y_width => 3
    )
    port map (
      x => delay1_q_net_x0,
      y => x3lsb_3_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/CRC Byte En/Skip First 2"

entity skip_first_2_entity_0ccfc7a7f5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    tx_reset: in std_logic; 
    en_2: out std_logic
  );
end skip_first_2_entity_0ccfc7a7f5;

architecture structural of skip_first_2_entity_0ccfc7a7f5 is
  signal ce_1_sg_x11: std_logic;
  signal clk_1_sg_x11: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x6: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;

begin
  ce_1_sg_x11 <= ce_1;
  clk_1_sg_x11 <= clk_1;
  logical1_y_net_x2 <= en;
  logical_y_net_x6 <= tx_reset;
  en_2 <= logical2_y_net_x0;

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x2,
      d1(0) => register2_q_net_x0,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x2,
      d1(0) => register2_q_net_x1,
      y(0) => logical2_y_net_x0
    );

  s_r_latch1_2f09b88201: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      r => logical_y_net_x6,
      s => logical1_y_net_x1,
      q => register2_q_net_x1
    );

  s_r_latch_6792cd308a: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x11,
      clk_1 => clk_1_sg_x11,
      r => logical_y_net_x6,
      s => logical1_y_net_x2,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/CRC Byte En"

entity crc_byte_en_entity_1ec74857a5 is
  port (
    bit_sel: in std_logic_vector(2 downto 0); 
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data: in std_logic; 
    logical_x0: in std_logic; 
    byte_en: out std_logic
  );
end crc_byte_en_entity_1ec74857a5;

architecture structural of crc_byte_en_entity_1ec74857a5 is
  signal ce_1_sg_x12: std_logic;
  signal clk_1_sg_x12: std_logic;
  signal constant3_op_net: std_logic_vector(1 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay_q_net_x0: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x7: std_logic;
  signal relational1_op_net: std_logic;
  signal x3lsb_y_net_x1: std_logic_vector(2 downto 0);

begin
  x3lsb_y_net_x1 <= bit_sel;
  delay_q_net_x0 <= bit_valid;
  ce_1_sg_x12 <= ce_1;
  clk_1_sg_x12 <= clk_1;
  delay2_q_net_x0 <= data;
  logical_y_net_x7 <= logical_x0;
  byte_en <= logical2_y_net_x1;

  constant3: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net_x0,
      d1(0) => delay_q_net_x0,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net,
      d1(0) => relational1_op_net,
      y(0) => logical1_y_net_x2
    );

  relational1: entity work.relational_632978e9ce
    port map (
      a => constant3_op_net,
      b => x3lsb_y_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  skip_first_2_0ccfc7a7f5: entity work.skip_first_2_entity_0ccfc7a7f5
    port map (
      ce_1 => ce_1_sg_x12,
      clk_1 => clk_1_sg_x12,
      en => logical1_y_net_x2,
      tx_reset => logical_y_net_x7,
      en_2 => logical2_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/CRC32 Calc/Endian Swap"

entity endian_swap_entity_227e3549f9 is
  port (
    b: in std_logic_vector(7 downto 0); 
    i: out std_logic_vector(7 downto 0)
  );
end endian_swap_entity_227e3549f9;

architecture structural of endian_swap_entity_227e3549f9 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b4_y_net: std_logic;
  signal b5_y_net: std_logic;
  signal b6_y_net: std_logic;
  signal b7_y_net: std_logic;
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal mux_y_net_x5: std_logic_vector(7 downto 0);

begin
  mux_y_net_x5 <= b;
  i <= concat_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b3_y_net
    );

  b4: entity work.xlslice
    generic map (
      new_lsb => 4,
      new_msb => 4,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b4_y_net
    );

  b5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 5,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b5_y_net
    );

  b6: entity work.xlslice
    generic map (
      new_lsb => 6,
      new_msb => 6,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b6_y_net
    );

  b7: entity work.xlslice
    generic map (
      new_lsb => 7,
      new_msb => 7,
      x_width => 8,
      y_width => 1
    )
    port map (
      x => mux_y_net_x5,
      y(0) => b7_y_net
    );

  concat: entity work.concat_7673b9b993
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => b0_y_net,
      in1(0) => b1_y_net,
      in2(0) => b2_y_net,
      in3(0) => b3_y_net,
      in4(0) => b4_y_net,
      in5(0) => b5_y_net,
      in6(0) => b6_y_net,
      in7(0) => b7_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b/CRC32 Calc"

entity crc32_calc_entity_7f133cdc7c is
  port (
    byte: in std_logic_vector(7 downto 0); 
    byte_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    tx_reset: in std_logic; 
    crc32: out std_logic_vector(31 downto 0)
  );
end crc32_calc_entity_7f133cdc7c;

architecture structural of crc32_calc_entity_7f133cdc7c is
  signal assert1_dout_net: std_logic_vector(31 downto 0);
  signal b0_y_net_x1: std_logic_vector(7 downto 0);
  signal b1_y_net_x1: std_logic_vector(7 downto 0);
  signal b2_y_net_x1: std_logic_vector(7 downto 0);
  signal b3_y_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x13: std_logic;
  signal clk_1_sg_x13: std_logic;
  signal concat1_y_net: std_logic_vector(31 downto 0);
  signal concat_y_net_x0: std_logic_vector(7 downto 0);
  signal concat_y_net_x1: std_logic_vector(7 downto 0);
  signal concat_y_net_x2: std_logic_vector(7 downto 0);
  signal concat_y_net_x3: std_logic_vector(7 downto 0);
  signal concat_y_net_x4: std_logic_vector(7 downto 0);
  signal concat_y_net_x5: std_logic_vector(31 downto 0);
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal crc_accum_q_net: std_logic_vector(31 downto 0);
  signal crc_remainders1_data_net: std_logic_vector(31 downto 0);
  signal inverter_op_net: std_logic_vector(31 downto 0);
  signal logical2_y_net_x2: std_logic;
  signal logical3_y_net: std_logic_vector(7 downto 0);
  signal logical4_y_net: std_logic_vector(31 downto 0);
  signal logical_y_net_x8: std_logic;
  signal mux_y_net_x6: std_logic_vector(7 downto 0);
  signal x24lsb_y_net: std_logic_vector(23 downto 0);
  signal x8msb_y_net: std_logic_vector(7 downto 0);

begin
  mux_y_net_x6 <= byte;
  logical2_y_net_x2 <= byte_valid;
  ce_1_sg_x13 <= ce_1;
  clk_1_sg_x13 <= clk_1;
  logical_y_net_x8 <= tx_reset;
  crc32 <= concat_y_net_x5;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 32,
      dout_width => 32
    )
    port map (
      din => crc_accum_q_net,
      dout => assert1_dout_net
    );

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b0_y_net_x1
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b1_y_net_x1
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b2_y_net_x1
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => inverter_op_net,
      y => b3_y_net_x1
    );

  concat: entity work.concat_a1e126f11c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => concat_y_net_x1,
      in1 => concat_y_net_x2,
      in2 => concat_y_net_x3,
      in3 => concat_y_net_x4,
      y => concat_y_net_x5
    );

  concat1: entity work.concat_c048fbe4a5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => x24lsb_y_net,
      in1 => constant1_op_net,
      y => concat1_y_net
    );

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  crc_accum: entity work.xlregister
    generic map (
      d_width => 32,
      init_value => b"11111111111111111111111111111111"
    )
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      d => logical4_y_net,
      en(0) => logical2_y_net_x2,
      rst(0) => logical_y_net_x8,
      q => crc_accum_q_net
    );

  crc_remainders1: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 8,
      c_address_width => 8,
      c_width => 32,
      core_name0 => "dmg_72_134e91999cae8947",
      latency => 0
    )
    port map (
      addr => logical3_y_net,
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      en => "1",
      data => crc_remainders1_data_net
    );

  endian_swap1_b278182efc: entity work.endian_swap_entity_227e3549f9
    port map (
      b => b0_y_net_x1,
      i => concat_y_net_x1
    );

  endian_swap2_a6b2c0f9fc: entity work.endian_swap_entity_227e3549f9
    port map (
      b => b1_y_net_x1,
      i => concat_y_net_x2
    );

  endian_swap3_4735cd3a69: entity work.endian_swap_entity_227e3549f9
    port map (
      b => b2_y_net_x1,
      i => concat_y_net_x3
    );

  endian_swap4_1f580e79cd: entity work.endian_swap_entity_227e3549f9
    port map (
      b => b3_y_net_x1,
      i => concat_y_net_x4
    );

  endian_swap_227e3549f9: entity work.endian_swap_entity_227e3549f9
    port map (
      b => mux_y_net_x6,
      i => concat_y_net_x0
    );

  inverter: entity work.inverter_6a3d3dd4e5
    port map (
      ce => ce_1_sg_x13,
      clk => clk_1_sg_x13,
      clr => '0',
      ip => assert1_dout_net,
      op => inverter_op_net
    );

  logical3: entity work.logical_59f8d33339
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => x8msb_y_net,
      d1 => concat_y_net_x0,
      y => logical3_y_net
    );

  logical4: entity work.logical_b23aa74086
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat1_y_net,
      d1 => crc_remainders1_data_net,
      y => logical4_y_net
    );

  x24lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 23,
      x_width => 32,
      y_width => 24
    )
    port map (
      x => assert1_dout_net,
      y => x24lsb_y_net
    );

  x8msb: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 31,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => assert1_dout_net,
      y => x8msb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Data Sel 64b"

entity data_sel_64b_entity_23f62948bd is
  port (
    bit_ind: in std_logic_vector(14 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data: in std_logic; 
    fcs: in std_logic; 
    logical: in std_logic; 
    pad_tail: in std_logic; 
    ram_64b: in std_logic_vector(63 downto 0); 
    ram_valid: in std_logic; 
    b: out std_logic
  );
end data_sel_64b_entity_23f62948bd;

architecture structural of data_sel_64b_entity_23f62948bd is
  signal assert_dout_net: std_logic_vector(31 downto 0);
  signal ce_1_sg_x14: std_logic;
  signal clk_1_sg_x14: std_logic;
  signal concat_y_net_x0: std_logic_vector(1 downto 0);
  signal concat_y_net_x5: std_logic_vector(31 downto 0);
  signal constant1_op_net: std_logic_vector(31 downto 0);
  signal delay1_q_net_x1: std_logic_vector(14 downto 0);
  signal delay2_q_net_x1: std_logic;
  signal delay5_q_net_x0: std_logic;
  signal delay_q_net_x1: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical_y_net_x9: std_logic;
  signal mux_y_net_x3: std_logic_vector(2 downto 0);
  signal mux_y_net_x4: std_logic;
  signal mux_y_net_x6: std_logic_vector(7 downto 0);
  signal mux_y_net_x7: std_logic_vector(63 downto 0);
  signal simulation_multiplexer_dout_net_x1: std_logic_vector(63 downto 0);
  signal x3lsb_y_net_x1: std_logic_vector(2 downto 0);

begin
  delay1_q_net_x1 <= bit_ind;
  ce_1_sg_x14 <= ce_1;
  clk_1_sg_x14 <= clk_1;
  delay2_q_net_x1 <= data;
  delay5_q_net_x0 <= fcs;
  logical_y_net_x9 <= logical;
  logical3_y_net_x0 <= pad_tail;
  simulation_multiplexer_dout_net_x1 <= ram_64b;
  delay_q_net_x1 <= ram_valid;
  b <= mux_y_net_x4;

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 32,
      dout_width => 32
    )
    port map (
      din => concat_y_net_x5,
      dout => assert_dout_net
    );

  bit_sel_2c3a4baaeb: entity work.bit_sel_entity_2c3a4baaeb
    port map (
      b => mux_y_net_x6,
      b_sel => x3lsb_y_net_x1,
      b_x0 => mux_y_net_x4
    );

  byte_sel_1b5e475260: entity work.byte_sel_entity_1b5e475260
    port map (
      b_sel => mux_y_net_x3,
      x64b => mux_y_net_x7,
      b => mux_y_net_x6
    );

  byte_sel_3a45df7438: entity work.byte_sel_entity_3a45df7438
    port map (
      bit_ind => delay1_q_net_x1,
      ce_1 => ce_1_sg_x14,
      clk_1 => clk_1_sg_x14,
      src_sel => concat_y_net_x0,
      tx_reset => logical_y_net_x9,
      sel => mux_y_net_x3
    );

  concat: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => logical3_y_net_x0,
      in1(0) => delay5_q_net_x0,
      y => concat_y_net_x0
    );

  constant1: entity work.constant_37567836aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  crc32_calc_7f133cdc7c: entity work.crc32_calc_entity_7f133cdc7c
    port map (
      byte => mux_y_net_x6,
      byte_valid => logical2_y_net_x2,
      ce_1 => ce_1_sg_x14,
      clk_1 => clk_1_sg_x14,
      tx_reset => logical_y_net_x9,
      crc32 => concat_y_net_x5
    );

  crc_byte_en_1ec74857a5: entity work.crc_byte_en_entity_1ec74857a5
    port map (
      bit_sel => x3lsb_y_net_x1,
      bit_valid => delay_q_net_x1,
      ce_1 => ce_1_sg_x14,
      clk_1 => clk_1_sg_x14,
      data => delay2_q_net_x1,
      logical_x0 => logical_y_net_x9,
      byte_en => logical2_y_net_x2
    );

  mux: entity work.mux_f3924dc817
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => simulation_multiplexer_dout_net_x1,
      d1 => assert_dout_net,
      d2 => constant1_op_net,
      sel => concat_y_net_x0,
      y => mux_y_net_x7
    );

  x3lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 15,
      y_width => 3
    )
    port map (
      x => delay1_q_net_x1,
      y => x3lsb_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/SIGNAL Capture/SIGNAL Slice/Endian Swap4"

entity endian_swap4_entity_9b5503b9d6 is
  port (
    b: in std_logic_vector(3 downto 0); 
    i: out std_logic_vector(3 downto 0)
  );
end endian_swap4_entity_9b5503b9d6;

architecture structural of endian_swap4_entity_9b5503b9d6 is
  signal b0_y_net: std_logic;
  signal b1_y_net: std_logic;
  signal b2_y_net: std_logic;
  signal b3_y_net: std_logic;
  signal b_3_0_y_net: std_logic_vector(3 downto 0);
  signal concat_y_net_x0: std_logic_vector(3 downto 0);

begin
  b_3_0_y_net <= b;
  i <= concat_y_net_x0;

  b0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => b_3_0_y_net,
      y(0) => b0_y_net
    );

  b1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => b_3_0_y_net,
      y(0) => b1_y_net
    );

  b2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => b_3_0_y_net,
      y(0) => b2_y_net
    );

  b3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 4,
      y_width => 1
    )
    port map (
      x => b_3_0_y_net,
      y(0) => b3_y_net
    );

  concat: entity work.concat_a0c7cd7a34
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => b0_y_net,
      in1(0) => b1_y_net,
      in2(0) => b2_y_net,
      in3(0) => b3_y_net,
      y => concat_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/SIGNAL Capture/SIGNAL Slice"

entity signal_slice_entity_a23045745d is
  port (
    s: in std_logic_vector(23 downto 0); 
    invalid: out std_logic; 
    length: out std_logic_vector(11 downto 0); 
    rate: out std_logic_vector(3 downto 0)
  );
end signal_slice_entity_a23045745d;

architecture structural of signal_slice_entity_a23045745d is
  signal b_16_5_y_net_x0: std_logic_vector(11 downto 0);
  signal b_23_18_y_net: std_logic_vector(5 downto 0);
  signal b_3_0_y_net: std_logic_vector(3 downto 0);
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal logical5_y_net_x0: std_logic;
  signal relational1_op_net: std_logic;
  signal relational2_op_net: std_logic;
  signal signal_q_net_x0: std_logic_vector(23 downto 0);

begin
  signal_q_net_x0 <= s;
  invalid <= logical5_y_net_x0;
  length <= b_16_5_y_net_x0;
  rate <= concat_y_net_x1;

  b_16_5: entity work.xlslice
    generic map (
      new_lsb => 5,
      new_msb => 16,
      x_width => 24,
      y_width => 12
    )
    port map (
      x => signal_q_net_x0,
      y => b_16_5_y_net_x0
    );

  b_23_18: entity work.xlslice
    generic map (
      new_lsb => 18,
      new_msb => 23,
      x_width => 24,
      y_width => 6
    )
    port map (
      x => signal_q_net_x0,
      y => b_23_18_y_net
    );

  b_3_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 24,
      y_width => 4
    )
    port map (
      x => signal_q_net_x0,
      y => b_3_0_y_net
    );

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_d6e645765a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  endian_swap4_9b5503b9d6: entity work.endian_swap4_entity_9b5503b9d6
    port map (
      b => b_3_0_y_net,
      i => concat_y_net_x1
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational2_op_net,
      d1(0) => relational1_op_net,
      y(0) => logical5_y_net_x0
    );

  relational1: entity work.relational_c49d820dc8
    port map (
      a => b_23_18_y_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  relational2: entity work.relational_43590be5cb
    port map (
      a => b_16_5_y_net_x0,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/SIGNAL Capture"

entity signal_capture_entity_4d07ad26ca is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data: in std_logic_vector(63 downto 0); 
    en: in std_logic; 
    tx_reset: in std_logic; 
    data_n_cbps: out std_logic_vector(8 downto 0); 
    data_n_dbps: out std_logic_vector(8 downto 0); 
    error: out std_logic; 
    signal_code_rate: out std_logic_vector(1 downto 0); 
    signal_length: out std_logic_vector(11 downto 0); 
    signal_mod_sel: out std_logic_vector(1 downto 0)
  );
end signal_capture_entity_4d07ad26ca;

architecture structural of signal_capture_entity_4d07ad26ca is
  signal b_16_5_y_net_x1: std_logic_vector(11 downto 0);
  signal b_2_1_y_net: std_logic_vector(1 downto 0);
  signal ce_1_sg_x18: std_logic;
  signal clk_1_sg_x18: std_logic;
  signal concat_y_net_x1: std_logic_vector(3 downto 0);
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic_vector(8 downto 0);
  signal convert3_dout_net_x1: std_logic_vector(8 downto 0);
  signal convert4_dout_net: std_logic;
  signal convert5_dout_net: std_logic;
  signal convert6_dout_net_x0: std_logic_vector(1 downto 0);
  signal convert_dout_net: std_logic_vector(3 downto 0);
  signal delay1_q_net: std_logic;
  signal delay3_q_net_x1: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x10: std_logic;
  signal mcode_code_rate_net: std_logic_vector(1 downto 0);
  signal mcode_mod_order_net: std_logic_vector(2 downto 0);
  signal mcode_n_cbps_net: std_logic_vector(8 downto 0);
  signal mcode_n_dbps_net: std_logic_vector(7 downto 0);
  signal mcode_valid_net: std_logic;
  signal register_q_net_x0: std_logic;
  signal signal_q_net_x0: std_logic_vector(23 downto 0);
  signal simulation_multiplexer_dout_net_x2: std_logic_vector(63 downto 0);
  signal x24lsb_y_net: std_logic_vector(23 downto 0);

begin
  ce_1_sg_x18 <= ce_1;
  clk_1_sg_x18 <= clk_1;
  simulation_multiplexer_dout_net_x2 <= data;
  delay3_q_net_x1 <= en;
  logical_y_net_x10 <= tx_reset;
  data_n_cbps <= convert2_dout_net_x0;
  data_n_dbps <= convert3_dout_net_x1;
  error <= register_q_net_x0;
  signal_code_rate <= convert6_dout_net_x0;
  signal_length <= b_16_5_y_net_x1;
  signal_mod_sel <= b_2_1_y_net;

  b_2_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 2,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => convert_dout_net,
      y => b_2_1_y_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 3,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 4,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din => mcode_mod_order_net,
      en => "1",
      dout => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din(0) => mcode_valid_net,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 9,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 9,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din => mcode_n_cbps_net,
      en => "1",
      dout => convert2_dout_net_x0
    );

  convert3: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 8,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 9,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din => mcode_n_dbps_net,
      en => "1",
      dout => convert3_dout_net_x1
    );

  convert4: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din(0) => logical_y_net_x10,
      en => "1",
      dout(0) => convert4_dout_net
    );

  convert5: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din(0) => delay1_q_net,
      en => "1",
      dout(0) => convert5_dout_net
    );

  convert6: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 2,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 2,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      din => mcode_code_rate_net,
      en => "1",
      dout => convert6_dout_net_x0
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      d(0) => logical1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      clr => '0',
      ip(0) => convert1_dout_net,
      op(0) => inverter_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => logical5_y_net_x0,
      y(0) => logical_y_net
    );

  mcode: entity work.mcode_block_b45edf5eb5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      signal_rate => concat_y_net_x1,
      code_rate => mcode_code_rate_net,
      mod_order => mcode_mod_order_net,
      n_cbps => mcode_n_cbps_net,
      n_dbps => mcode_n_dbps_net,
      valid(0) => mcode_valid_net
    );

  posedge_c85fd78403: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x18,
      clk_1 => clk_1_sg_x18,
      d => delay3_q_net_x1,
      q => logical1_y_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      d(0) => logical_y_net,
      en(0) => convert5_dout_net,
      rst(0) => convert4_dout_net,
      q(0) => register_q_net_x0
    );

  signal_slice_a23045745d: entity work.signal_slice_entity_a23045745d
    port map (
      s => signal_q_net_x0,
      invalid => logical5_y_net_x0,
      length => b_16_5_y_net_x1,
      rate => concat_y_net_x1
    );

  signal_x0: entity work.xlregister
    generic map (
      d_width => 24,
      init_value => b"000000000001000000001010"
    )
    port map (
      ce => ce_1_sg_x18,
      clk => clk_1_sg_x18,
      d => x24lsb_y_net,
      en(0) => logical1_y_net_x0,
      rst(0) => logical_y_net_x10,
      q => signal_q_net_x0
    );

  x24lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 23,
      x_width => 64,
      y_width => 24
    )
    port map (
      x => simulation_multiplexer_dout_net_x2,
      y => x24lsb_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source/Sym Compute Ctrl"

entity sym_compute_ctrl_entity_03292a0793 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    last_bit_in_sym: in std_logic; 
    output_fifo_occ: in std_logic_vector(7 downto 0); 
    regtx_cp_len: in std_logic_vector(7 downto 0); 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    tx_iq_samp_ce: in std_logic; 
    tx_reset: in std_logic; 
    tx_running: in std_logic; 
    start_next_sym: out std_logic
  );
end sym_compute_ctrl_entity_03292a0793;

architecture structural of sym_compute_ctrl_entity_03292a0793 is
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal b_15_8_y_net: std_logic_vector(7 downto 0);
  signal b_7_0_y_net: std_logic_vector(7 downto 0);
  signal ce_1_sg_x24: std_logic;
  signal clk_1_sg_x24: std_logic;
  signal constant_op_net: std_logic_vector(7 downto 0);
  signal convert2_dout_net_x0: std_logic;
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal delay2_q_net: std_logic;
  signal fifo_dcount_net_x0: std_logic_vector(7 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal inverter_op_net_x3: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical6_y_net: std_logic;
  signal logical_y_net_x12: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x2: std_logic;
  signal register2_q_net_x3: std_logic;
  signal relational2_op_net_x0: std_logic;
  signal relational3_op_net: std_logic;

begin
  ce_1_sg_x24 <= ce_1;
  clk_1_sg_x24 <= clk_1;
  inverter_op_net_x3 <= last_bit_in_sym;
  fifo_dcount_net_x0 <= output_fifo_occ;
  b_15_8_y_net <= regtx_cp_len;
  b_7_0_y_net <= regtx_num_sc;
  convert2_dout_net_x0 <= tx_iq_samp_ce;
  logical_y_net_x12 <= tx_reset;
  register2_q_net_x3 <= tx_running;
  start_next_sym <= logical1_y_net_x4;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 8,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 9,
      core_name0 => "addsb_11_0_8dc9188fad4d9a9c",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 9,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => b_7_0_y_net,
      b => b_15_8_y_net,
      ce => ce_1_sg_x24,
      clk => clk_1_sg_x24,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant_x0: entity work.constant_c936744458
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_d24951bef2f0cdc9",
      op_arith => xlUnsigned,
      op_width => 7
    )
    port map (
      ce => ce_1_sg_x24,
      clk => clk_1_sg_x24,
      clr => '0',
      en(0) => logical4_y_net,
      rst(0) => logical6_y_net,
      op => counter_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 80,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x24,
      clk => clk_1_sg_x24,
      d(0) => logical2_y_net,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x24,
      clk => clk_1_sg_x24,
      clr => '0',
      ip(0) => register2_q_net_x0,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x24,
      clk => clk_1_sg_x24,
      clr => '0',
      ip(0) => register2_q_net_x3,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_a6d07705dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x0,
      d1(0) => delay2_q_net,
      d2(0) => logical3_y_net,
      d3(0) => logical1_y_net_x3,
      y(0) => logical1_y_net_x4
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net_x3,
      d1(0) => inverter_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => register2_q_net_x3,
      d2(0) => relational3_op_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x2,
      d1(0) => convert2_dout_net_x0,
      y(0) => logical4_y_net
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter1_op_net,
      d1(0) => logical_y_net_x12,
      y(0) => logical5_y_net_x0
    );

  logical6: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => logical_y_net_x12,
      y(0) => logical6_y_net
    );

  posedge1_92cf7422b9: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x24,
      clk_1 => clk_1_sg_x24,
      d => relational2_op_net_x0,
      q => logical1_y_net_x1
    );

  posedge2_215c090ff9: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x24,
      clk_1 => clk_1_sg_x24,
      d => register2_q_net_x2,
      q => logical1_y_net_x3
    );

  posedge_53b708e5e5: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x24,
      clk_1 => clk_1_sg_x24,
      d => register2_q_net_x3,
      q => logical1_y_net_x0
    );

  relational2: entity work.relational_5a9c998b07
    port map (
      a => fifo_dcount_net_x0,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net_x0
    );

  relational3: entity work.relational_19bf67ea71
    port map (
      a => counter_op_net,
      b => addsub_s_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_d224ea7cc5: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x24,
      clk_1 => clk_1_sg_x24,
      r => logical5_y_net_x0,
      s => logical1_y_net_x1,
      q => register2_q_net_x2
    );

  s_r_latch_d1eaca1541: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x24,
      clk_1 => clk_1_sg_x24,
      r => logical_y_net_x12,
      s => inverter_op_net_x3,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Bit Source"

entity bit_source_entity_8a38dc99ff is
  port (
    b_15_8: in std_logic_vector(7 downto 0); 
    b_23_16: in std_logic_vector(7 downto 0); 
    b_7_0: in std_logic_vector(7 downto 0); 
    bram_din: in std_logic_vector(63 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    convert2: in std_logic; 
    done: in std_logic; 
    fifo: in std_logic_vector(7 downto 0); 
    mux: in std_logic_vector(3 downto 0); 
    tx_reset: in std_logic; 
    tx_start: in std_logic; 
    addr_gen: out std_logic; 
    bit: out std_logic; 
    bit_valid: out std_logic; 
    bram_if_64b: out std_logic_vector(31 downto 0); 
    bram_if_64b_x0: out std_logic; 
    bram_if_64b_x1: out std_logic; 
    bram_if_64b_x2: out std_logic_vector(63 downto 0); 
    bram_if_64b_x3: out std_logic_vector(7 downto 0); 
    data_pad_fcs: out std_logic; 
    signal_capture: out std_logic_vector(8 downto 0); 
    signal_capture_x0: out std_logic_vector(1 downto 0); 
    signal_capture_x1: out std_logic_vector(1 downto 0); 
    signal_decode_error: out std_logic; 
    tail: out std_logic
  );
end bit_source_entity_8a38dc99ff;

architecture structural of bit_source_entity_8a38dc99ff is
  signal accumulator_q_net_x1: std_logic_vector(14 downto 0);
  signal b_15_8_y_net_x0: std_logic_vector(7 downto 0);
  signal b_16_5_y_net_x1: std_logic_vector(11 downto 0);
  signal b_23_16_y_net_x1: std_logic_vector(7 downto 0);
  signal b_2_1_y_net_x0: std_logic_vector(1 downto 0);
  signal b_7_0_y_net_x0: std_logic_vector(7 downto 0);
  signal bram_din_net_x1: std_logic_vector(63 downto 0);
  signal ce_1_sg_x25: std_logic;
  signal clk_1_sg_x25: std_logic;
  signal concat_y_net_x1: std_logic_vector(31 downto 0);
  signal constant1_op_net_x1: std_logic;
  signal constant2_op_net_x1: std_logic;
  signal constant7_op_net_x1: std_logic_vector(63 downto 0);
  signal constant8_op_net_x1: std_logic_vector(7 downto 0);
  signal convert2_dout_net_x2: std_logic;
  signal convert2_dout_net_x3: std_logic_vector(8 downto 0);
  signal convert3_dout_net_x1: std_logic_vector(8 downto 0);
  signal convert6_dout_net_x1: std_logic_vector(1 downto 0);
  signal delay1_q_net_x1: std_logic_vector(14 downto 0);
  signal delay2_q_net_x1: std_logic;
  signal delay3_q_net_x1: std_logic;
  signal delay3_q_net_x2: std_logic;
  signal delay3_q_net_x3: std_logic;
  signal delay4_q_net_x0: std_logic;
  signal delay5_q_net_x0: std_logic;
  signal delay6_q_net: std_logic;
  signal delay_q_net_x2: std_logic;
  signal fifo_dcount_net_x1: std_logic_vector(7 downto 0);
  signal inverter_op_net_x3: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal logical3_y_net_x1: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical_y_net_x1: std_logic;
  signal logical_y_net_x13: std_logic;
  signal mux_y_net_x1: std_logic_vector(3 downto 0);
  signal mux_y_net_x5: std_logic;
  signal register2_q_net_x3: std_logic;
  signal register_q_net_x1: std_logic;
  signal register_q_net_x2: std_logic;
  signal relational6_op_net_x0: std_logic;
  signal simulation_multiplexer_dout_net_x2: std_logic_vector(63 downto 0);

begin
  b_15_8_y_net_x0 <= b_15_8;
  b_23_16_y_net_x1 <= b_23_16;
  b_7_0_y_net_x0 <= b_7_0;
  bram_din_net_x1 <= bram_din;
  ce_1_sg_x25 <= ce_1;
  clk_1_sg_x25 <= clk_1;
  convert2_dout_net_x2 <= convert2;
  delay3_q_net_x2 <= done;
  fifo_dcount_net_x1 <= fifo;
  mux_y_net_x1 <= mux;
  logical_y_net_x13 <= tx_reset;
  logical_y_net_x1 <= tx_start;
  addr_gen <= delay3_q_net_x3;
  bit <= mux_y_net_x5;
  bit_valid <= delay_q_net_x2;
  bram_if_64b <= concat_y_net_x1;
  bram_if_64b_x0 <= constant1_op_net_x1;
  bram_if_64b_x1 <= constant2_op_net_x1;
  bram_if_64b_x2 <= constant7_op_net_x1;
  bram_if_64b_x3 <= constant8_op_net_x1;
  data_pad_fcs <= logical1_y_net_x2;
  signal_capture <= convert2_dout_net_x3;
  signal_capture_x0 <= convert6_dout_net_x1;
  signal_capture_x1 <= b_2_1_y_net_x0;
  signal_decode_error <= register_q_net_x1;
  tail <= delay4_q_net_x0;

  addr_gen_b968174b41: entity work.addr_gen_entity_b968174b41
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      en => register_q_net_x2,
      signal_length => b_16_5_y_net_x1,
      tx_reset => logical_y_net_x13,
      bit_mem_addr => accumulator_q_net_x1,
      data => logical2_y_net_x0,
      fcs => logical1_y_net_x0,
      pad => relational6_op_net_x0,
      ppdu_tail_done => delay3_q_net_x3,
      signal_x0 => logical5_y_net_x0,
      tail => logical3_y_net_x0
    );

  bit_per_sym_counter_be13008040: entity work.bit_per_sym_counter_entity_be13008040
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      data_n_dbps => convert3_dout_net_x1,
      start_sym => logical1_y_net_x4,
      tx_reset => logical_y_net_x13,
      last_bit_in_sym => inverter_op_net_x3,
      load_bit => register_q_net_x2
    );

  bram_if_64b_672a3af05d: entity work.bram_if_64b_entity_672a3af05d
    port map (
      bit_addr => accumulator_q_net_x1,
      bram_din => bram_din_net_x1,
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      regtx_pkt_buf_addr_offset => b_23_16_y_net_x1,
      tx_pkt_buf_sel => mux_y_net_x1,
      concat_x0 => concat_y_net_x1,
      constant1_x0 => constant1_op_net_x1,
      constant2_x0 => constant2_op_net_x1,
      constant7_x0 => constant7_op_net_x1,
      constant8_x0 => constant8_op_net_x1,
      x64b_data => simulation_multiplexer_dout_net_x2
    );

  data_sel_64b_23f62948bd: entity work.data_sel_64b_entity_23f62948bd
    port map (
      bit_ind => delay1_q_net_x1,
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      data => delay2_q_net_x1,
      fcs => delay5_q_net_x0,
      logical => logical_y_net_x13,
      pad_tail => logical3_y_net_x1,
      ram_64b => simulation_multiplexer_dout_net_x2,
      ram_valid => delay_q_net_x2,
      b => mux_y_net_x5
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => register_q_net_x2,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x2
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 15
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d => accumulator_q_net_x1,
      en => '1',
      rst => '1',
      q => delay1_q_net_x1
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => logical2_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x1
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => logical5_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x1
    );

  delay4: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => logical3_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay4_q_net_x0
    );

  delay5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => logical1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay5_q_net_x0
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x25,
      clk => clk_1_sg_x25,
      d(0) => relational6_op_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net
    );

  logical1: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net_x1,
      d1(0) => delay6_q_net,
      d2(0) => delay5_q_net_x0,
      y(0) => logical1_y_net_x2
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x13,
      d1(0) => delay3_q_net_x2,
      y(0) => logical2_y_net_x1
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay4_q_net_x0,
      d1(0) => delay6_q_net,
      y(0) => logical3_y_net_x1
    );

  posedge_8f9c4e7e37: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      d => logical_y_net_x1,
      q => logical1_y_net_x1
    );

  s_r_latch_4263c9ab1a: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      r => logical2_y_net_x1,
      s => logical1_y_net_x1,
      q => register2_q_net_x3
    );

  signal_capture_4d07ad26ca: entity work.signal_capture_entity_4d07ad26ca
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      data => simulation_multiplexer_dout_net_x2,
      en => delay3_q_net_x1,
      tx_reset => logical_y_net_x13,
      data_n_cbps => convert2_dout_net_x3,
      data_n_dbps => convert3_dout_net_x1,
      error => register_q_net_x1,
      signal_code_rate => convert6_dout_net_x1,
      signal_length => b_16_5_y_net_x1,
      signal_mod_sel => b_2_1_y_net_x0
    );

  sym_compute_ctrl_03292a0793: entity work.sym_compute_ctrl_entity_03292a0793
    port map (
      ce_1 => ce_1_sg_x25,
      clk_1 => clk_1_sg_x25,
      last_bit_in_sym => inverter_op_net_x3,
      output_fifo_occ => fifo_dcount_net_x1,
      regtx_cp_len => b_15_8_y_net_x0,
      regtx_num_sc => b_7_0_y_net_x0,
      tx_iq_samp_ce => convert2_dout_net_x2,
      tx_reset => logical_y_net_x13,
      tx_running => register2_q_net_x3,
      start_next_sym => logical1_y_net_x4
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/EDK Processor"

entity edk_processor_entity_de00edcbbe is
  port (
    axi_aresetn: in std_logic; 
    from_register: in std_logic_vector(31 downto 0); 
    plb_ce_1: in std_logic; 
    plb_clk_1: in std_logic; 
    s_axi_araddr: in std_logic_vector(31 downto 0); 
    s_axi_arburst: in std_logic_vector(1 downto 0); 
    s_axi_arcache: in std_logic_vector(3 downto 0); 
    s_axi_arid: in std_logic_vector(7 downto 0); 
    s_axi_arlen: in std_logic_vector(7 downto 0); 
    s_axi_arlock: in std_logic_vector(1 downto 0); 
    s_axi_arprot: in std_logic_vector(2 downto 0); 
    s_axi_arsize: in std_logic_vector(2 downto 0); 
    s_axi_arvalid: in std_logic; 
    s_axi_awaddr: in std_logic_vector(31 downto 0); 
    s_axi_awburst: in std_logic_vector(1 downto 0); 
    s_axi_awcache: in std_logic_vector(3 downto 0); 
    s_axi_awid: in std_logic_vector(7 downto 0); 
    s_axi_awlen: in std_logic_vector(7 downto 0); 
    s_axi_awlock: in std_logic_vector(1 downto 0); 
    s_axi_awprot: in std_logic_vector(2 downto 0); 
    s_axi_awsize: in std_logic_vector(2 downto 0); 
    s_axi_awvalid: in std_logic; 
    s_axi_bready: in std_logic; 
    s_axi_rready: in std_logic; 
    s_axi_wdata: in std_logic_vector(31 downto 0); 
    s_axi_wlast: in std_logic; 
    s_axi_wstrb: in std_logic_vector(3 downto 0); 
    s_axi_wvalid: in std_logic; 
    to_register: in std_logic_vector(31 downto 0); 
    to_register1: in std_logic_vector(31 downto 0); 
    to_register2: in std_logic_vector(31 downto 0); 
    to_register3: in std_logic_vector(31 downto 0); 
    to_register4: in std_logic_vector(31 downto 0); 
    to_register5: in std_logic_vector(31 downto 0); 
    memmap_x0: out std_logic; 
    memmap_x1: out std_logic; 
    memmap_x10: out std_logic; 
    memmap_x11: out std_logic_vector(31 downto 0); 
    memmap_x12: out std_logic; 
    memmap_x13: out std_logic_vector(31 downto 0); 
    memmap_x14: out std_logic; 
    memmap_x15: out std_logic_vector(31 downto 0); 
    memmap_x16: out std_logic; 
    memmap_x17: out std_logic_vector(31 downto 0); 
    memmap_x18: out std_logic; 
    memmap_x19: out std_logic_vector(31 downto 0); 
    memmap_x2: out std_logic_vector(7 downto 0); 
    memmap_x20: out std_logic; 
    memmap_x21: out std_logic_vector(31 downto 0); 
    memmap_x22: out std_logic; 
    memmap_x3: out std_logic_vector(1 downto 0); 
    memmap_x4: out std_logic; 
    memmap_x5: out std_logic_vector(31 downto 0); 
    memmap_x6: out std_logic_vector(7 downto 0); 
    memmap_x7: out std_logic; 
    memmap_x8: out std_logic_vector(1 downto 0); 
    memmap_x9: out std_logic
  );
end edk_processor_entity_de00edcbbe;

architecture structural of edk_processor_entity_de00edcbbe is
  signal axi_aresetn_net_x0: std_logic;
  signal from_register_data_out_net_x0: std_logic_vector(31 downto 0);
  signal memmap_s_axi_arready_net_x0: std_logic;
  signal memmap_s_axi_awready_net_x0: std_logic;
  signal memmap_s_axi_bid_net_x0: std_logic_vector(7 downto 0);
  signal memmap_s_axi_bresp_net_x0: std_logic_vector(1 downto 0);
  signal memmap_s_axi_bvalid_net_x0: std_logic;
  signal memmap_s_axi_rdata_net_x0: std_logic_vector(31 downto 0);
  signal memmap_s_axi_rid_net_x0: std_logic_vector(7 downto 0);
  signal memmap_s_axi_rlast_net_x0: std_logic;
  signal memmap_s_axi_rresp_net_x0: std_logic_vector(1 downto 0);
  signal memmap_s_axi_rvalid_net_x0: std_logic;
  signal memmap_s_axi_wready_net_x0: std_logic;
  signal memmap_sm_config_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_config_en_net_x0: std_logic;
  signal memmap_sm_fft_config_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_fft_config_en_net_x0: std_logic;
  signal memmap_sm_output_scaling_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_output_scaling_en_net_x0: std_logic;
  signal memmap_sm_pkt_buf_sel_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_pkt_buf_sel_en_net_x0: std_logic;
  signal memmap_sm_timing_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_timing_en_net_x0: std_logic;
  signal memmap_sm_tx_start_din_net_x0: std_logic_vector(31 downto 0);
  signal memmap_sm_tx_start_en_net_x0: std_logic;
  signal plb_ce_1_sg_x0: std_logic;
  signal plb_clk_1_sg_x0: std_logic;
  signal s_axi_araddr_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_arburst_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_arcache_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_arid_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_arlen_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_arlock_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_arprot_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_arsize_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_arvalid_net_x0: std_logic;
  signal s_axi_awaddr_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_awburst_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_awcache_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_awid_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_awlen_net_x0: std_logic_vector(7 downto 0);
  signal s_axi_awlock_net_x0: std_logic_vector(1 downto 0);
  signal s_axi_awprot_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_awsize_net_x0: std_logic_vector(2 downto 0);
  signal s_axi_awvalid_net_x0: std_logic;
  signal s_axi_bready_net_x0: std_logic;
  signal s_axi_rready_net_x0: std_logic;
  signal s_axi_wdata_net_x0: std_logic_vector(31 downto 0);
  signal s_axi_wlast_net_x0: std_logic;
  signal s_axi_wstrb_net_x0: std_logic_vector(3 downto 0);
  signal s_axi_wvalid_net_x0: std_logic;
  signal to_register1_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register2_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register3_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register4_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register5_dout_net_x0: std_logic_vector(31 downto 0);
  signal to_register_dout_net_x0: std_logic_vector(31 downto 0);

begin
  axi_aresetn_net_x0 <= axi_aresetn;
  from_register_data_out_net_x0 <= from_register;
  plb_ce_1_sg_x0 <= plb_ce_1;
  plb_clk_1_sg_x0 <= plb_clk_1;
  s_axi_araddr_net_x0 <= s_axi_araddr;
  s_axi_arburst_net_x0 <= s_axi_arburst;
  s_axi_arcache_net_x0 <= s_axi_arcache;
  s_axi_arid_net_x0 <= s_axi_arid;
  s_axi_arlen_net_x0 <= s_axi_arlen;
  s_axi_arlock_net_x0 <= s_axi_arlock;
  s_axi_arprot_net_x0 <= s_axi_arprot;
  s_axi_arsize_net_x0 <= s_axi_arsize;
  s_axi_arvalid_net_x0 <= s_axi_arvalid;
  s_axi_awaddr_net_x0 <= s_axi_awaddr;
  s_axi_awburst_net_x0 <= s_axi_awburst;
  s_axi_awcache_net_x0 <= s_axi_awcache;
  s_axi_awid_net_x0 <= s_axi_awid;
  s_axi_awlen_net_x0 <= s_axi_awlen;
  s_axi_awlock_net_x0 <= s_axi_awlock;
  s_axi_awprot_net_x0 <= s_axi_awprot;
  s_axi_awsize_net_x0 <= s_axi_awsize;
  s_axi_awvalid_net_x0 <= s_axi_awvalid;
  s_axi_bready_net_x0 <= s_axi_bready;
  s_axi_rready_net_x0 <= s_axi_rready;
  s_axi_wdata_net_x0 <= s_axi_wdata;
  s_axi_wlast_net_x0 <= s_axi_wlast;
  s_axi_wstrb_net_x0 <= s_axi_wstrb;
  s_axi_wvalid_net_x0 <= s_axi_wvalid;
  to_register_dout_net_x0 <= to_register;
  to_register1_dout_net_x0 <= to_register1;
  to_register2_dout_net_x0 <= to_register2;
  to_register3_dout_net_x0 <= to_register3;
  to_register4_dout_net_x0 <= to_register4;
  to_register5_dout_net_x0 <= to_register5;
  memmap_x0 <= memmap_s_axi_arready_net_x0;
  memmap_x1 <= memmap_s_axi_awready_net_x0;
  memmap_x10 <= memmap_s_axi_wready_net_x0;
  memmap_x11 <= memmap_sm_timing_din_net_x0;
  memmap_x12 <= memmap_sm_timing_en_net_x0;
  memmap_x13 <= memmap_sm_config_din_net_x0;
  memmap_x14 <= memmap_sm_config_en_net_x0;
  memmap_x15 <= memmap_sm_pkt_buf_sel_din_net_x0;
  memmap_x16 <= memmap_sm_pkt_buf_sel_en_net_x0;
  memmap_x17 <= memmap_sm_output_scaling_din_net_x0;
  memmap_x18 <= memmap_sm_output_scaling_en_net_x0;
  memmap_x19 <= memmap_sm_tx_start_din_net_x0;
  memmap_x2 <= memmap_s_axi_bid_net_x0;
  memmap_x20 <= memmap_sm_tx_start_en_net_x0;
  memmap_x21 <= memmap_sm_fft_config_din_net_x0;
  memmap_x22 <= memmap_sm_fft_config_en_net_x0;
  memmap_x3 <= memmap_s_axi_bresp_net_x0;
  memmap_x4 <= memmap_s_axi_bvalid_net_x0;
  memmap_x5 <= memmap_s_axi_rdata_net_x0;
  memmap_x6 <= memmap_s_axi_rid_net_x0;
  memmap_x7 <= memmap_s_axi_rlast_net_x0;
  memmap_x8 <= memmap_s_axi_rresp_net_x0;
  memmap_x9 <= memmap_s_axi_rvalid_net_x0;

  memmap: entity work.axi_sgiface
    port map (
      axi_aclk => plb_clk_1_sg_x0,
      axi_aresetn => axi_aresetn_net_x0,
      axi_ce => plb_ce_1_sg_x0,
      s_axi_araddr => s_axi_araddr_net_x0,
      s_axi_arburst => s_axi_arburst_net_x0,
      s_axi_arcache => s_axi_arcache_net_x0,
      s_axi_arid => s_axi_arid_net_x0,
      s_axi_arlen => s_axi_arlen_net_x0,
      s_axi_arlock => s_axi_arlock_net_x0,
      s_axi_arprot => s_axi_arprot_net_x0,
      s_axi_arsize => s_axi_arsize_net_x0,
      s_axi_arvalid => s_axi_arvalid_net_x0,
      s_axi_awaddr => s_axi_awaddr_net_x0,
      s_axi_awburst => s_axi_awburst_net_x0,
      s_axi_awcache => s_axi_awcache_net_x0,
      s_axi_awid => s_axi_awid_net_x0,
      s_axi_awlen => s_axi_awlen_net_x0,
      s_axi_awlock => s_axi_awlock_net_x0,
      s_axi_awprot => s_axi_awprot_net_x0,
      s_axi_awsize => s_axi_awsize_net_x0,
      s_axi_awvalid => s_axi_awvalid_net_x0,
      s_axi_bready => s_axi_bready_net_x0,
      s_axi_rready => s_axi_rready_net_x0,
      s_axi_wdata => s_axi_wdata_net_x0,
      s_axi_wlast => s_axi_wlast_net_x0,
      s_axi_wstrb => s_axi_wstrb_net_x0,
      s_axi_wvalid => s_axi_wvalid_net_x0,
      sm_config_dout => to_register1_dout_net_x0,
      sm_fft_config_dout => to_register5_dout_net_x0,
      sm_output_scaling_dout => to_register3_dout_net_x0,
      sm_pkt_buf_sel_dout => to_register2_dout_net_x0,
      sm_status_dout => from_register_data_out_net_x0,
      sm_timing_dout => to_register_dout_net_x0,
      sm_tx_start_dout => to_register4_dout_net_x0,
      s_axi_arready => memmap_s_axi_arready_net_x0,
      s_axi_awready => memmap_s_axi_awready_net_x0,
      s_axi_bid => memmap_s_axi_bid_net_x0,
      s_axi_bresp => memmap_s_axi_bresp_net_x0,
      s_axi_bvalid => memmap_s_axi_bvalid_net_x0,
      s_axi_rdata => memmap_s_axi_rdata_net_x0,
      s_axi_rid => memmap_s_axi_rid_net_x0,
      s_axi_rlast => memmap_s_axi_rlast_net_x0,
      s_axi_rresp => memmap_s_axi_rresp_net_x0,
      s_axi_rvalid => memmap_s_axi_rvalid_net_x0,
      s_axi_wready => memmap_s_axi_wready_net_x0,
      sm_config_din => memmap_sm_config_din_net_x0,
      sm_config_en => memmap_sm_config_en_net_x0,
      sm_fft_config_din => memmap_sm_fft_config_din_net_x0,
      sm_fft_config_en => memmap_sm_fft_config_en_net_x0,
      sm_output_scaling_din => memmap_sm_output_scaling_din_net_x0,
      sm_output_scaling_en => memmap_sm_output_scaling_en_net_x0,
      sm_pkt_buf_sel_din => memmap_sm_pkt_buf_sel_din_net_x0,
      sm_pkt_buf_sel_en => memmap_sm_pkt_buf_sel_en_net_x0,
      sm_timing_din => memmap_sm_timing_din_net_x0,
      sm_timing_en => memmap_sm_timing_en_net_x0,
      sm_tx_start_din => memmap_sm_tx_start_din_net_x0,
      sm_tx_start_en => memmap_sm_tx_start_en_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/FFT/FFT Core"

entity fft_core_entity_0a10ef78f5 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_in_tlast: in std_logic; 
    data_in_tvalid: in std_logic; 
    i_in: in std_logic_vector(15 downto 0); 
    q_in: in std_logic_vector(15 downto 0); 
    regtx_cp_len: in std_logic_vector(7 downto 0); 
    regtx_fft_scaling: in std_logic_vector(5 downto 0); 
    tx_reset: in std_logic; 
    data_in_tready: out std_logic; 
    data_out_tlast: out std_logic; 
    data_out_tvalid: out std_logic; 
    i_out: out std_logic_vector(15 downto 0); 
    q_out: out std_logic_vector(15 downto 0)
  );
end fft_core_entity_0a10ef78f5;

architecture structural of fft_core_entity_0a10ef78f5 is
  signal axi_fifo_m_axis_tvalid_net_x0: std_logic;
  signal b_15_8_y_net_x1: std_logic_vector(7 downto 0);
  signal b_29_24_y_net: std_logic_vector(5 downto 0);
  signal ce_1_sg_x26: std_logic;
  signal clk_1_sg_x26: std_logic;
  signal constant1_op_net: std_logic;
  signal constant2_op_net: std_logic;
  signal constant3_op_net: std_logic;
  signal constant4_op_net: std_logic;
  signal convert_dout_net: std_logic_vector(5 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x0: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x0: std_logic;
  signal inverter_op_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x14: std_logic;
  signal reinterpret2_output_port_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x0: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x26 <= ce_1;
  clk_1_sg_x26 <= clk_1;
  logical2_y_net_x0 <= data_in_tlast;
  axi_fifo_m_axis_tvalid_net_x0 <= data_in_tvalid;
  reinterpret2_output_port_net_x0 <= i_in;
  reinterpret3_output_port_net_x0 <= q_in;
  b_15_8_y_net_x1 <= regtx_cp_len;
  b_29_24_y_net <= regtx_fft_scaling;
  logical_y_net_x14 <= tx_reset;
  data_in_tready <= fast_fourier_transform_8_0_s_axis_data_tready_net_x0;
  data_out_tlast <= fast_fourier_transform_8_0_m_axis_data_tlast_net_x0;
  data_out_tvalid <= fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0;
  i_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0;
  q_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0;

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant2: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  constant3: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant3_op_net
    );

  constant4: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant4_op_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 8,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 6,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x26,
      clk => clk_1_sg_x26,
      clr => '0',
      din => b_15_8_y_net_x1,
      en => "1",
      dout => convert_dout_net
    );

  fast_fourier_transform_8_0: entity work.xlfast_fourier_transform_66965782653510ded5a0002b36532651
    port map (
      ce => ce_1_sg_x26,
      clk => clk_1_sg_x26,
      m_axis_data_tready => constant3_op_net,
      m_axis_status_tready => constant2_op_net,
      rst => inverter_op_net,
      s_axis_config_tdata_cp_len => convert_dout_net,
      s_axis_config_tdata_fwd_inv(0) => constant1_op_net,
      s_axis_config_tdata_scale_sch => b_29_24_y_net,
      s_axis_config_tvalid => constant4_op_net,
      s_axis_data_tdata_xn_im => reinterpret3_output_port_net_x0,
      s_axis_data_tdata_xn_re => reinterpret2_output_port_net_x0,
      s_axis_data_tlast => logical2_y_net_x0,
      s_axis_data_tvalid => axi_fifo_m_axis_tvalid_net_x0,
      m_axis_data_tdata_xk_im => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x0,
      m_axis_data_tdata_xk_re => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x0,
      m_axis_data_tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x0,
      m_axis_data_tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x0,
      s_axis_data_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x0
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x26,
      clk => clk_1_sg_x26,
      clr => '0',
      ip(0) => logical_y_net_x14,
      op(0) => inverter_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/FFT"

entity fft_entity_b2c6e5af27 is
  port (
    b_15_8: in std_logic_vector(7 downto 0); 
    b_29_24: in std_logic_vector(5 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_in_tlast: in std_logic; 
    data_in_tvalid: in std_logic; 
    i_in: in std_logic_vector(15 downto 0); 
    last_sym: in std_logic; 
    q_in: in std_logic_vector(15 downto 0); 
    tx_reset: in std_logic; 
    data_in_tready: out std_logic; 
    data_out_tvalid: out std_logic; 
    i_out: out std_logic_vector(15 downto 0); 
    last_sym_x0: out std_logic; 
    q_out: out std_logic_vector(15 downto 0)
  );
end fft_entity_b2c6e5af27;

architecture structural of fft_entity_b2c6e5af27 is
  signal axi_fifo_m_axis_tvalid_net_x1: std_logic;
  signal b_15_8_y_net_x2: std_logic_vector(7 downto 0);
  signal b_29_24_y_net_x0: std_logic_vector(5 downto 0);
  signal ce_1_sg_x28: std_logic;
  signal clk_1_sg_x28: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tlast_net_x0: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x1: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x16: std_logic;
  signal register2_q_net_x0: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(15 downto 0);

begin
  b_15_8_y_net_x2 <= b_15_8;
  b_29_24_y_net_x0 <= b_29_24;
  ce_1_sg_x28 <= ce_1;
  clk_1_sg_x28 <= clk_1;
  logical2_y_net_x1 <= data_in_tlast;
  axi_fifo_m_axis_tvalid_net_x1 <= data_in_tvalid;
  reinterpret2_output_port_net_x1 <= i_in;
  logical1_y_net_x1 <= last_sym;
  reinterpret3_output_port_net_x1 <= q_in;
  logical_y_net_x16 <= tx_reset;
  data_in_tready <= fast_fourier_transform_8_0_s_axis_data_tready_net_x1;
  data_out_tvalid <= fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1;
  i_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1;
  last_sym_x0 <= logical_y_net_x0;
  q_out <= fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1;

  fft_core_0a10ef78f5: entity work.fft_core_entity_0a10ef78f5
    port map (
      ce_1 => ce_1_sg_x28,
      clk_1 => clk_1_sg_x28,
      data_in_tlast => logical2_y_net_x1,
      data_in_tvalid => axi_fifo_m_axis_tvalid_net_x1,
      i_in => reinterpret2_output_port_net_x1,
      q_in => reinterpret3_output_port_net_x1,
      regtx_cp_len => b_15_8_y_net_x2,
      regtx_fft_scaling => b_29_24_y_net_x0,
      tx_reset => logical_y_net_x16,
      data_in_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x1,
      data_out_tlast => fast_fourier_transform_8_0_m_axis_data_tlast_net_x0,
      data_out_tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x1,
      i_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x1,
      q_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x1
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => fast_fourier_transform_8_0_m_axis_data_tlast_net_x0,
      d1(0) => register2_q_net_x0,
      y(0) => logical_y_net_x0
    );

  s_r_latch2_ec8501d2e6: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x28,
      clk_1 => clk_1_sg_x28,
      r => logical_y_net_x16,
      s => logical1_y_net_x1,
      q => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/FIFO/I/Q Concat"

entity q_concat_entity_e63daf7dbb is
  port (
    i: in std_logic_vector(15 downto 0); 
    q: in std_logic_vector(15 downto 0); 
    iq: out std_logic_vector(31 downto 0)
  );
end q_concat_entity_e63daf7dbb;

architecture structural of q_concat_entity_e63daf7dbb is
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert1_dout_net_x0: std_logic_vector(15 downto 0);
  signal convert_dout_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  convert_dout_net_x0 <= i;
  convert1_dout_net_x0 <= q;
  iq <= concat_y_net_x0;

  concat: entity work.concat_a369e00c6b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net_x0
    );

  reinterpret: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_dout_net_x0,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert1_dout_net_x0,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/FIFO/I/Q Slice"

entity q_slice_entity_10657a6c34 is
  port (
    iq: in std_logic_vector(31 downto 0); 
    i: out std_logic_vector(15 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end q_slice_entity_10657a6c34;

architecture structural of q_slice_entity_10657a6c34 is
  signal axi_fifo_m_axis_tdata_net_x0: std_logic_vector(31 downto 0);
  signal reinterpret2_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x2: std_logic_vector(15 downto 0);
  signal slice1_y_net: std_logic_vector(15 downto 0);
  signal slice_y_net: std_logic_vector(15 downto 0);

begin
  axi_fifo_m_axis_tdata_net_x0 <= iq;
  i <= reinterpret2_output_port_net_x2;
  q <= reinterpret3_output_port_net_x2;

  reinterpret2: entity work.reinterpret_151459306d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice_y_net,
      output_port => reinterpret2_output_port_net_x2
    );

  reinterpret3: entity work.reinterpret_151459306d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => slice1_y_net,
      output_port => reinterpret3_output_port_net_x2
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 31,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => axi_fifo_m_axis_tdata_net_x0,
      y => slice_y_net
    );

  slice1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 15,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => axi_fifo_m_axis_tdata_net_x0,
      y => slice1_y_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/FIFO"

entity fifo_entity_c992f1a4af is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_tvalid: in std_logic; 
    fft_tready: in std_logic; 
    i: in std_logic_vector(11 downto 0); 
    last_samp: in std_logic; 
    last_sym: in std_logic; 
    q: in std_logic_vector(11 downto 0); 
    tx_reset: in std_logic; 
    fft_tdata_im: out std_logic_vector(15 downto 0); 
    fft_tdata_re: out std_logic_vector(15 downto 0); 
    fft_tlast: out std_logic; 
    fft_tvalid: out std_logic; 
    fifo_tready: out std_logic; 
    last_sym_x0: out std_logic
  );
end fifo_entity_c992f1a4af;

architecture structural of fifo_entity_c992f1a4af is
  signal axi_fifo_m_axis_tdata_net_x0: std_logic_vector(31 downto 0);
  signal axi_fifo_m_axis_tlast_net: std_logic;
  signal axi_fifo_m_axis_tuser_net: std_logic;
  signal axi_fifo_m_axis_tvalid_net_x2: std_logic;
  signal axi_fifo_s_axis_tready_net_x0: std_logic;
  signal ce_1_sg_x29: std_logic;
  signal clk_1_sg_x29: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert1_dout_net_x0: std_logic_vector(15 downto 0);
  signal convert2_dout_net: std_logic;
  signal convert3_dout_net: std_logic;
  signal convert_dout_net_x0: std_logic_vector(15 downto 0);
  signal delay1_q_net_x0: std_logic;
  signal delay3_q_net_x3: std_logic;
  signal delay_q_net_x0: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x2: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal logical_y_net_x17: std_logic;
  signal mux3_y_net_x0: std_logic_vector(11 downto 0);
  signal mux4_y_net_x0: std_logic_vector(11 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x3: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x29 <= ce_1;
  clk_1_sg_x29 <= clk_1;
  delay_q_net_x0 <= data_tvalid;
  fast_fourier_transform_8_0_s_axis_data_tready_net_x2 <= fft_tready;
  mux3_y_net_x0 <= i;
  delay1_q_net_x0 <= last_samp;
  delay3_q_net_x3 <= last_sym;
  mux4_y_net_x0 <= q;
  logical_y_net_x17 <= tx_reset;
  fft_tdata_im <= reinterpret3_output_port_net_x3;
  fft_tdata_re <= reinterpret2_output_port_net_x3;
  fft_tlast <= logical2_y_net_x2;
  fft_tvalid <= axi_fifo_m_axis_tvalid_net_x2;
  fifo_tready <= axi_fifo_s_axis_tready_net_x0;
  last_sym_x0 <= logical1_y_net_x2;

  axi_fifo: entity work.xlaxififogen_wlan_phy_tx_pmd
    generic map (
      core_name0 => "axififo_fg92_4d50ffea04713b7c",
      depth_bits => 7,
      has_aresetn => 1,
      tdata_width => 32,
      tuser_width => 1
    )
    port map (
      aresetn => inverter_op_net,
      ce => ce_1_sg_x29,
      m_axis_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x2,
      s_aclk => clk_1_sg_x29,
      s_axis_tdata => concat_y_net_x0,
      s_axis_tlast => delay1_q_net_x0,
      s_axis_tuser(0) => convert2_dout_net,
      s_axis_tvalid => delay_q_net_x0,
      m_axis_tdata => axi_fifo_m_axis_tdata_net_x0,
      m_axis_tlast => axi_fifo_m_axis_tlast_net,
      m_axis_tuser(0) => axi_fifo_m_axis_tuser_net,
      m_axis_tvalid => axi_fifo_m_axis_tvalid_net_x2,
      s_axis_tready => axi_fifo_s_axis_tready_net_x0
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 11,
      din_width => 12,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din => mux3_y_net_x0,
      en => "1",
      dout => convert_dout_net_x0
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 11,
      din_width => 12,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din => mux4_y_net_x0,
      en => "1",
      dout => convert1_dout_net_x0
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din(0) => delay3_q_net_x3,
      en => "1",
      dout(0) => convert2_dout_net
    );

  convert3: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      din(0) => axi_fifo_m_axis_tuser_net,
      en => "1",
      dout(0) => convert3_dout_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x29,
      clk => clk_1_sg_x29,
      clr => '0',
      ip(0) => logical_y_net_x17,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => axi_fifo_m_axis_tvalid_net_x2,
      d1(0) => convert3_dout_net,
      y(0) => logical1_y_net_x2
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => axi_fifo_m_axis_tvalid_net_x2,
      d1(0) => axi_fifo_m_axis_tlast_net,
      y(0) => logical2_y_net_x2
    );

  q_concat_e63daf7dbb: entity work.q_concat_entity_e63daf7dbb
    port map (
      i => convert_dout_net_x0,
      q => convert1_dout_net_x0,
      iq => concat_y_net_x0
    );

  q_slice_10657a6c34: entity work.q_slice_entity_10657a6c34
    port map (
      iq => axi_fifo_m_axis_tdata_net_x0,
      i => reinterpret2_output_port_net_x3,
      q => reinterpret3_output_port_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/16-QAM/16QAM Int Addr/Osc"

entity osc_entity_4b2508a4db is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    r: in std_logic; 
    q: out std_logic
  );
end osc_entity_4b2508a4db;

architecture structural of osc_entity_4b2508a4db is
  signal assert_dout_net: std_logic;
  signal ce_1_sg_x30: std_logic;
  signal clk_1_sg_x30: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical_y_net_x18: std_logic;
  signal register2_q_net_x0: std_logic;

begin
  ce_1_sg_x30 <= ce_1;
  clk_1_sg_x30 <= clk_1;
  logical1_y_net_x0 <= en;
  logical_y_net_x18 <= r;
  q <= register2_q_net_x0;

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register2_q_net_x0,
      dout(0) => assert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      din(0) => logical_y_net_x18,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      din(0) => logical1_y_net_x0,
      en => "1",
      dout(0) => convert2_dout_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      clr => '0',
      ip(0) => assert_dout_net,
      op(0) => inverter_op_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x30,
      clk => clk_1_sg_x30,
      d(0) => inverter_op_net,
      en(0) => convert2_dout_net,
      rst(0) => convert1_dout_net,
      q(0) => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/16-QAM/16QAM Int Addr"

entity x16qam_int_addr_entity_f990691d0d is
  port (
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    new_sym: in std_logic; 
    tx_reset: in std_logic; 
    wr_addr: out std_logic_vector(7 downto 0); 
    wr_offset: out std_logic
  );
end x16qam_int_addr_entity_f990691d0d;

architecture structural of x16qam_int_addr_entity_f990691d0d is
  signal ce_1_sg_x32: std_logic;
  signal clk_1_sg_x32: std_logic;
  signal constant2_op_net: std_logic_vector(7 downto 0);
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal delay2_q_net_x1: std_logic;
  signal delay2_q_net_x2: std_logic;
  signal delay_q_net_x0: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x19: std_logic;
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;
  signal x16qam_ind_data_net_x0: std_logic_vector(7 downto 0);

begin
  delay_q_net_x0 <= bit_valid;
  ce_1_sg_x32 <= ce_1;
  clk_1_sg_x32 <= clk_1;
  delay2_q_net_x1 <= new_sym;
  logical_y_net_x19 <= tx_reset;
  wr_addr <= x16qam_ind_data_net_x0;
  wr_offset <= delay2_q_net_x2;

  constant2: entity work.constant_6e2bcf24f9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 191,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_86806e294f737f4c",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      clr => '0',
      en(0) => delay_q_net_x0,
      rst(0) => logical1_y_net,
      op => counter_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x2
    );

  logical1: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x19,
      d1(0) => delay2_q_net_x1,
      d2(0) => logical1_y_net_x1,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x0,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  osc_4b2508a4db: entity work.osc_entity_4b2508a4db
    port map (
      ce_1 => ce_1_sg_x32,
      clk_1 => clk_1_sg_x32,
      en => logical1_y_net_x1,
      r => logical_y_net_x19,
      q => register2_q_net_x0
    );

  posedge_a817475926: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x32,
      clk_1 => clk_1_sg_x32,
      d => logical2_y_net_x0,
      q => logical1_y_net_x1
    );

  relational2: entity work.relational_54048c8b02
    port map (
      a => counter_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  x16qam_ind: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 8,
      c_width => 8,
      core_name0 => "bmg_72_28f68c2bb9b4d938",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x32,
      clk => clk_1_sg_x32,
      en => "1",
      rst => "0",
      data => x16qam_ind_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/16-QAM"

entity x16_qam_entity_381a479990 is
  port (
    bit_tdata: in std_logic; 
    bit_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_sym_addr: in std_logic_vector(5 downto 0); 
    logical: in std_logic; 
    new_sym: in std_logic; 
    x4b_data: out std_logic_vector(3 downto 0)
  );
end x16_qam_entity_381a479990;

architecture structural of x16_qam_entity_381a479990 is
  signal bit_memory1_doutb_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x33: std_logic;
  signal clk_1_sg_x33: std_logic;
  signal concat1_y_net: std_logic_vector(8 downto 0);
  signal concat2_y_net: std_logic_vector(6 downto 0);
  signal constant1_op_net: std_logic_vector(3 downto 0);
  signal constant2_op_net: std_logic;
  signal delay2_q_net: std_logic;
  signal delay2_q_net_x2: std_logic;
  signal delay2_q_net_x3: std_logic;
  signal delay6_q_net: std_logic;
  signal delay_q_net_x1: std_logic;
  signal inverter_op_net: std_logic;
  signal logical_y_net_x20: std_logic;
  signal mux_y_net_x0: std_logic;
  signal slice_y_net_x0: std_logic_vector(5 downto 0);
  signal x16qam_ind_data_net_x0: std_logic_vector(7 downto 0);

begin
  mux_y_net_x0 <= bit_tdata;
  delay_q_net_x1 <= bit_tvalid;
  ce_1_sg_x33 <= ce_1;
  clk_1_sg_x33 <= clk_1;
  slice_y_net_x0 <= data_sym_addr;
  logical_y_net_x20 <= logical;
  delay2_q_net_x3 <= new_sym;
  x4b_data <= bit_memory1_doutb_net_x0;

  bit_memory1: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 9,
      c_address_width_b => 7,
      c_width_a => 1,
      c_width_b => 4,
      core_name0 => "bmg_72_7ec9033b751d2879",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x33,
      a_clk => clk_1_sg_x33,
      addra => concat1_y_net,
      addrb => concat2_y_net,
      b_ce => ce_1_sg_x33,
      b_clk => clk_1_sg_x33,
      dina(0) => delay6_q_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => delay2_q_net,
      web(0) => constant2_op_net,
      doutb => bit_memory1_doutb_net_x0
    );

  concat1: entity work.concat_1ece14600f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay2_q_net_x2,
      in1 => x16qam_ind_data_net_x0,
      y => concat1_y_net
    );

  concat2: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => inverter_op_net,
      in1 => slice_y_net_x0,
      y => concat2_y_net
    );

  constant1: entity work.constant_4c449dd556
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      d(0) => delay_q_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      d(0) => mux_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x33,
      clk => clk_1_sg_x33,
      clr => '0',
      ip(0) => delay2_q_net_x2,
      op(0) => inverter_op_net
    );

  x16qam_int_addr_f990691d0d: entity work.x16qam_int_addr_entity_f990691d0d
    port map (
      bit_valid => delay_q_net_x1,
      ce_1 => ce_1_sg_x33,
      clk_1 => clk_1_sg_x33,
      new_sym => delay2_q_net_x3,
      tx_reset => logical_y_net_x20,
      wr_addr => x16qam_ind_data_net_x0,
      wr_offset => delay2_q_net_x2
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/16QAM Mod"

entity x16qam_mod_entity_cce570a88c is
  port (
    b_3_0: in std_logic_vector(3 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end x16qam_mod_entity_cce570a88c;

architecture structural of x16qam_mod_entity_cce570a88c is
  signal b_1_0_y_net: std_logic_vector(1 downto 0);
  signal b_3_2_y_net: std_logic_vector(1 downto 0);
  signal bit_memory1_doutb_net_x1: std_logic_vector(3 downto 0);
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);

begin
  bit_memory1_doutb_net_x1 <= b_3_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  b_1_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 1,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => bit_memory1_doutb_net_x1,
      y => b_1_0_y_net
    );

  b_3_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 3,
      x_width => 4,
      y_width => 2
    )
    port map (
      x => bit_memory1_doutb_net_x1,
      y => b_3_2_y_net
    );

  constant1: entity work.constant_8cac5f7cf5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_1bebc71bf9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_92715f6857
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_9b9cbaee60
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  mux: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      sel => b_1_0_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      sel => b_3_2_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/64-QAM/64QAM Int Addr"

entity x64qam_int_addr_entity_dcc862cdc9 is
  port (
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    new_sym: in std_logic; 
    tx_reset: in std_logic; 
    wr_addr: out std_logic_vector(8 downto 0); 
    wr_offset: out std_logic
  );
end x64qam_int_addr_entity_dcc862cdc9;

architecture structural of x64qam_int_addr_entity_dcc862cdc9 is
  signal ce_1_sg_x36: std_logic;
  signal clk_1_sg_x36: std_logic;
  signal constant2_op_net: std_logic_vector(8 downto 0);
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x4: std_logic;
  signal delay_q_net_x2: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x22: std_logic;
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;
  signal x64qam_ind_data_net_x0: std_logic_vector(8 downto 0);

begin
  delay_q_net_x2 <= bit_valid;
  ce_1_sg_x36 <= ce_1;
  clk_1_sg_x36 <= clk_1;
  delay2_q_net_x4 <= new_sym;
  logical_y_net_x22 <= tx_reset;
  wr_addr <= x64qam_ind_data_net_x0;
  wr_offset <= delay2_q_net_x0;

  constant2: entity work.constant_8d143efc5e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 287,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_36e2bb554c95560d",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      clr => '0',
      en(0) => delay_q_net_x2,
      rst(0) => logical1_y_net,
      op => counter_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  logical1: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x22,
      d1(0) => delay2_q_net_x4,
      d2(0) => logical1_y_net_x1,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x2,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  osc_edab26a8af: entity work.osc_entity_4b2508a4db
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      en => logical1_y_net_x1,
      r => logical_y_net_x22,
      q => register2_q_net_x0
    );

  posedge_8bc118b07b: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x36,
      clk_1 => clk_1_sg_x36,
      d => logical2_y_net_x0,
      q => logical1_y_net_x1
    );

  relational2: entity work.relational_6c3ee657fa
    port map (
      a => counter_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  x64qam_ind: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 9,
      c_width => 9,
      core_name0 => "bmg_72_324b883165919716",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x36,
      clk => clk_1_sg_x36,
      en => "1",
      rst => "0",
      data => x64qam_ind_data_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/64-QAM"

entity x64_qam_entity_35dea913c2 is
  port (
    bit_tdata: in std_logic; 
    bit_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_sym_addr: in std_logic_vector(5 downto 0); 
    logical: in std_logic; 
    new_sym: in std_logic; 
    x6b_data: out std_logic_vector(5 downto 0)
  );
end x64_qam_entity_35dea913c2;

architecture structural of x64_qam_entity_35dea913c2 is
  signal bit_memory1_doutb_net: std_logic_vector(7 downto 0);
  signal ce_1_sg_x37: std_logic;
  signal clk_1_sg_x37: std_logic;
  signal concat1_y_net: std_logic_vector(9 downto 0);
  signal concat2_y_net: std_logic_vector(6 downto 0);
  signal constant1_op_net: std_logic_vector(7 downto 0);
  signal constant2_op_net: std_logic;
  signal delay2_q_net: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x5: std_logic;
  signal delay6_q_net: std_logic;
  signal delay_q_net_x3: std_logic;
  signal inverter_op_net: std_logic;
  signal logical_y_net_x23: std_logic;
  signal mux_y_net_x1: std_logic;
  signal slice_y_net_x1: std_logic_vector(5 downto 0);
  signal slice_y_net_x2: std_logic_vector(5 downto 0);
  signal x64qam_ind_data_net_x0: std_logic_vector(8 downto 0);

begin
  mux_y_net_x1 <= bit_tdata;
  delay_q_net_x3 <= bit_tvalid;
  ce_1_sg_x37 <= ce_1;
  clk_1_sg_x37 <= clk_1;
  slice_y_net_x1 <= data_sym_addr;
  logical_y_net_x23 <= logical;
  delay2_q_net_x5 <= new_sym;
  x6b_data <= slice_y_net_x2;

  bit_memory1: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 10,
      c_address_width_b => 7,
      c_width_a => 1,
      c_width_b => 8,
      core_name0 => "bmg_72_da153342fc52049b",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x37,
      a_clk => clk_1_sg_x37,
      addra => concat1_y_net,
      addrb => concat2_y_net,
      b_ce => ce_1_sg_x37,
      b_clk => clk_1_sg_x37,
      dina(0) => delay6_q_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => delay2_q_net,
      web(0) => constant2_op_net,
      doutb => bit_memory1_doutb_net
    );

  concat1: entity work.concat_9779a5cf83
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay2_q_net_x0,
      in1 => x64qam_ind_data_net_x0,
      y => concat1_y_net
    );

  concat2: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => inverter_op_net,
      in1 => slice_y_net_x1,
      y => concat2_y_net
    );

  constant1: entity work.constant_91ef1678ca
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      d(0) => delay_q_net_x3,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      d(0) => mux_y_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x37,
      clk => clk_1_sg_x37,
      clr => '0',
      ip(0) => delay2_q_net_x0,
      op(0) => inverter_op_net
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 8,
      y_width => 6
    )
    port map (
      x => bit_memory1_doutb_net,
      y => slice_y_net_x2
    );

  x64qam_int_addr_dcc862cdc9: entity work.x64qam_int_addr_entity_dcc862cdc9
    port map (
      bit_valid => delay_q_net_x3,
      ce_1 => ce_1_sg_x37,
      clk_1 => clk_1_sg_x37,
      new_sym => delay2_q_net_x5,
      tx_reset => logical_y_net_x23,
      wr_addr => x64qam_ind_data_net_x0,
      wr_offset => delay2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/64QAM Mod"

entity x64qam_mod_entity_e734ca01a6 is
  port (
    b_5_0: in std_logic_vector(5 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end x64qam_mod_entity_e734ca01a6;

architecture structural of x64qam_mod_entity_e734ca01a6 is
  signal b_2_0_y_net: std_logic_vector(2 downto 0);
  signal b_5_3_y_net: std_logic_vector(2 downto 0);
  signal constant10_op_net: std_logic_vector(11 downto 0);
  signal constant11_op_net: std_logic_vector(11 downto 0);
  signal constant12_op_net: std_logic_vector(11 downto 0);
  signal constant13_op_net: std_logic_vector(11 downto 0);
  signal constant14_op_net: std_logic_vector(11 downto 0);
  signal constant15_op_net: std_logic_vector(11 downto 0);
  signal constant16_op_net: std_logic_vector(11 downto 0);
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net: std_logic_vector(11 downto 0);
  signal constant5_op_net: std_logic_vector(11 downto 0);
  signal constant6_op_net: std_logic_vector(11 downto 0);
  signal constant7_op_net: std_logic_vector(11 downto 0);
  signal constant8_op_net: std_logic_vector(11 downto 0);
  signal constant9_op_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal slice_y_net_x3: std_logic_vector(5 downto 0);

begin
  slice_y_net_x3 <= b_5_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  b_2_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 2,
      x_width => 6,
      y_width => 3
    )
    port map (
      x => slice_y_net_x3,
      y => b_2_0_y_net
    );

  b_5_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 5,
      x_width => 6,
      y_width => 3
    )
    port map (
      x => slice_y_net_x3,
      y => b_5_3_y_net
    );

  constant1: entity work.constant_9127ce6619
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant10: entity work.constant_555e35158a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant10_op_net
    );

  constant11: entity work.constant_c0e78ca39c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant11_op_net
    );

  constant12: entity work.constant_e3898a7c17
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant12_op_net
    );

  constant13: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant13_op_net
    );

  constant14: entity work.constant_d3e8ce78bb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant14_op_net
    );

  constant15: entity work.constant_20bb1d9cec
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant15_op_net
    );

  constant16: entity work.constant_044e9822dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant16_op_net
    );

  constant2: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_d3e8ce78bb
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_20bb1d9cec
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  constant5: entity work.constant_9127ce6619
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_555e35158a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  constant7: entity work.constant_c0e78ca39c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant7_op_net
    );

  constant8: entity work.constant_e3898a7c17
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant8_op_net
    );

  constant9: entity work.constant_044e9822dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant9_op_net
    );

  mux: entity work.mux_f3bb14635d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant1_op_net,
      d2 => constant3_op_net,
      d3 => constant4_op_net,
      d4 => constant10_op_net,
      d5 => constant9_op_net,
      d6 => constant11_op_net,
      d7 => constant12_op_net,
      sel => b_2_0_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_f3bb14635d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant13_op_net,
      d1 => constant5_op_net,
      d2 => constant14_op_net,
      d3 => constant15_op_net,
      d4 => constant6_op_net,
      d5 => constant16_op_net,
      d6 => constant7_op_net,
      d7 => constant8_op_net,
      sel => b_5_3_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/BPSK/BPSK Int Addr"

entity bpsk_int_addr_entity_c4e932a6e5 is
  port (
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    new_sym: in std_logic; 
    tx_reset: in std_logic; 
    wr_addr: out std_logic_vector(5 downto 0); 
    wr_offset: out std_logic
  );
end bpsk_int_addr_entity_c4e932a6e5;

architecture structural of bpsk_int_addr_entity_c4e932a6e5 is
  signal bpsk_int_data_net_x0: std_logic_vector(5 downto 0);
  signal ce_1_sg_x40: std_logic;
  signal clk_1_sg_x40: std_logic;
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal counter_op_net: std_logic_vector(5 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x6: std_logic;
  signal delay_q_net_x4: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x25: std_logic;
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;

begin
  delay_q_net_x4 <= bit_valid;
  ce_1_sg_x40 <= ce_1;
  clk_1_sg_x40 <= clk_1;
  delay2_q_net_x6 <= new_sym;
  logical_y_net_x25 <= tx_reset;
  wr_addr <= bpsk_int_data_net_x0;
  wr_offset <= delay2_q_net_x0;

  bpsk_int: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 6,
      c_width => 6,
      core_name0 => "bmg_72_f580ae3be5511d30",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      en => "1",
      rst => "0",
      data => bpsk_int_data_net_x0
    );

  constant2: entity work.constant_ef95fb0eb4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 47,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_f068fb73312ae1e5",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      clr => '0',
      en(0) => delay_q_net_x4,
      rst(0) => logical1_y_net,
      op => counter_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x40,
      clk => clk_1_sg_x40,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  logical1: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x25,
      d1(0) => delay2_q_net_x6,
      d2(0) => logical1_y_net_x1,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x4,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  osc_f7a0ec6b9b: entity work.osc_entity_4b2508a4db
    port map (
      ce_1 => ce_1_sg_x40,
      clk_1 => clk_1_sg_x40,
      en => logical1_y_net_x1,
      r => logical_y_net_x25,
      q => register2_q_net_x0
    );

  posedge_7e7b4014a8: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x40,
      clk_1 => clk_1_sg_x40,
      d => logical2_y_net_x0,
      q => logical1_y_net_x1
    );

  relational2: entity work.relational_931d61fb72
    port map (
      a => counter_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/BPSK"

entity bpsk_entity_ba0b27afd0 is
  port (
    bit_tdata: in std_logic; 
    bit_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_sym_addr: in std_logic_vector(5 downto 0); 
    logical: in std_logic; 
    new_sym: in std_logic; 
    x1b_data: out std_logic
  );
end bpsk_entity_ba0b27afd0;

architecture structural of bpsk_entity_ba0b27afd0 is
  signal bit_memory_doutb_net_x0: std_logic;
  signal bpsk_int_data_net_x0: std_logic_vector(5 downto 0);
  signal ce_1_sg_x41: std_logic;
  signal clk_1_sg_x41: std_logic;
  signal concat1_y_net: std_logic_vector(6 downto 0);
  signal concat2_y_net: std_logic_vector(6 downto 0);
  signal constant1_op_net: std_logic;
  signal constant2_op_net: std_logic;
  signal delay1_q_net: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x7: std_logic;
  signal delay6_q_net: std_logic;
  signal delay_q_net_x5: std_logic;
  signal inverter_op_net: std_logic;
  signal logical_y_net_x26: std_logic;
  signal mux_y_net_x2: std_logic;
  signal slice_y_net_x2: std_logic_vector(5 downto 0);

begin
  mux_y_net_x2 <= bit_tdata;
  delay_q_net_x5 <= bit_tvalid;
  ce_1_sg_x41 <= ce_1;
  clk_1_sg_x41 <= clk_1;
  slice_y_net_x2 <= data_sym_addr;
  logical_y_net_x26 <= logical;
  delay2_q_net_x7 <= new_sym;
  x1b_data <= bit_memory_doutb_net_x0;

  bit_memory: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 7,
      c_address_width_b => 7,
      c_width_a => 1,
      c_width_b => 1,
      core_name0 => "bmg_72_41985f385eaacb3e",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x41,
      a_clk => clk_1_sg_x41,
      addra => concat1_y_net,
      addrb => concat2_y_net,
      b_ce => ce_1_sg_x41,
      b_clk => clk_1_sg_x41,
      dina(0) => delay6_q_net,
      dinb(0) => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => delay1_q_net,
      web(0) => constant2_op_net,
      doutb(0) => bit_memory_doutb_net_x0
    );

  bpsk_int_addr_c4e932a6e5: entity work.bpsk_int_addr_entity_c4e932a6e5
    port map (
      bit_valid => delay_q_net_x5,
      ce_1 => ce_1_sg_x41,
      clk_1 => clk_1_sg_x41,
      new_sym => delay2_q_net_x7,
      tx_reset => logical_y_net_x26,
      wr_addr => bpsk_int_data_net_x0,
      wr_offset => delay2_q_net_x0
    );

  concat1: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay2_q_net_x0,
      in1 => bpsk_int_data_net_x0,
      y => concat1_y_net
    );

  concat2: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => inverter_op_net,
      in1 => slice_y_net_x2,
      y => concat2_y_net
    );

  constant1: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      d(0) => delay_q_net_x5,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      d(0) => mux_y_net_x2,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x41,
      clk => clk_1_sg_x41,
      clr => '0',
      ip(0) => delay2_q_net_x0,
      op(0) => inverter_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/BPSK Mod"

entity bpsk_mod_entity_9dd399b8d9 is
  port (
    b_0: in std_logic; 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end bpsk_mod_entity_9dd399b8d9;

architecture structural of bpsk_mod_entity_9dd399b8d9 is
  signal bit_memory_doutb_net_x1: std_logic;
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal constant4_op_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);

begin
  bit_memory_doutb_net_x1 <= b_0;
  i <= mux_y_net_x0;
  q <= constant4_op_net_x0;

  constant2: entity work.constant_58c7454693
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_504d9a75aa
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net_x0
    );

  mux: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => bit_memory_doutb_net_x1,
      y => mux_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Coded Bit Counter"

entity coded_bit_counter_entity_bb3901367b is
  port (
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_n_cbps: in std_logic_vector(8 downto 0); 
    tx_reset: in std_logic; 
    bits_ready: out std_logic
  );
end coded_bit_counter_entity_bb3901367b;

architecture structural of coded_bit_counter_entity_bb3901367b is
  signal ce_1_sg_x43: std_logic;
  signal clk_1_sg_x43: std_logic;
  signal constant3_op_net: std_logic_vector(5 downto 0);
  signal convert2_dout_net_x4: std_logic_vector(8 downto 0);
  signal delay2_q_net_x8: std_logic;
  signal delay_q_net_x6: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x28: std_logic;
  signal mux_y_net: std_logic_vector(8 downto 0);
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;
  signal sym_coded_bit_count_op_net: std_logic_vector(8 downto 0);

begin
  delay_q_net_x6 <= bit_valid;
  ce_1_sg_x43 <= ce_1;
  clk_1_sg_x43 <= clk_1;
  convert2_dout_net_x4 <= data_n_cbps;
  logical_y_net_x28 <= tx_reset;
  bits_ready <= delay2_q_net_x8;

  constant3: entity work.constant_5c27e02321
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      d(0) => logical2_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x8
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      ip(0) => relational2_op_net,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical2_y_net_x0,
      d1(0) => logical_y_net_x28,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter_op_net,
      d1(0) => delay_q_net_x6,
      y(0) => logical2_y_net_x0
    );

  mux: entity work.mux_4075671a27
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant3_op_net,
      d1 => convert2_dout_net_x4,
      sel(0) => register2_q_net_x0,
      y => mux_y_net
    );

  relational2: entity work.relational_82fb466a8b
    port map (
      a => sym_coded_bit_count_op_net,
      b => mux_y_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  s_r_latch2_562a909877: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x43,
      clk_1 => clk_1_sg_x43,
      r => logical_y_net_x28,
      s => logical2_y_net_x0,
      q => register2_q_net_x0
    );

  sym_coded_bit_count: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_d66925a45384983e",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x43,
      clk => clk_1_sg_x43,
      clr => '0',
      en(0) => delay_q_net_x6,
      rst(0) => logical1_y_net,
      op => sym_coded_bit_count_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots/Data SC Map"

entity data_sc_map_entity_0f52ca1546 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    sc_ind: in std_logic_vector(5 downto 0); 
    data_sym_ind: out std_logic_vector(5 downto 0); 
    data_sym_valid: out std_logic
  );
end data_sc_map_entity_0f52ca1546;

architecture structural of data_sc_map_entity_0f52ca1546 is
  signal ce_1_sg_x44: std_logic;
  signal clk_1_sg_x44: std_logic;
  signal constant2_op_net: std_logic_vector(6 downto 0);
  signal relational1_op_net_x0: std_logic;
  signal sc_sym_map_data_net: std_logic_vector(6 downto 0);
  signal slice_y_net_x3: std_logic_vector(5 downto 0);
  signal subcarrier_index_op_net_x0: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x44 <= ce_1;
  clk_1_sg_x44 <= clk_1;
  subcarrier_index_op_net_x0 <= sc_ind;
  data_sym_ind <= slice_y_net_x3;
  data_sym_valid <= relational1_op_net_x0;

  constant2: entity work.constant_7b07120b87
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  relational1: entity work.relational_23065a6aa3
    port map (
      a => constant2_op_net,
      b => sc_sym_map_data_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  sc_sym_map: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 6,
      c_address_width => 6,
      c_width => 7,
      core_name0 => "dmg_72_5efcdb43c0011b51",
      latency => 0
    )
    port map (
      addr => subcarrier_index_op_net_x0,
      ce => ce_1_sg_x44,
      clk => clk_1_sg_x44,
      en => "1",
      data => sc_sym_map_data_net
    );

  slice: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 5,
      x_width => 7,
      y_width => 6
    )
    port map (
      x => sc_sym_map_data_net,
      y => slice_y_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots/Pilot Gen/Pilot Selection"

entity pilot_selection_entity_93fec99adc is
  port (
    sc_ind: in std_logic_vector(5 downto 0); 
    negate: out std_logic; 
    pilot: out std_logic
  );
end pilot_selection_entity_93fec99adc;

architecture structural of pilot_selection_entity_93fec99adc is
  signal constant1_op_net: std_logic_vector(5 downto 0);
  signal constant2_op_net: std_logic_vector(5 downto 0);
  signal constant3_op_net: std_logic_vector(5 downto 0);
  signal constant4_op_net: std_logic_vector(5 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal relational4_op_net: std_logic;
  signal relational5_op_net_x0: std_logic;
  signal relational6_op_net: std_logic;
  signal relational7_op_net: std_logic;
  signal subcarrier_index_op_net_x1: std_logic_vector(5 downto 0);

begin
  subcarrier_index_op_net_x1 <= sc_ind;
  negate <= relational5_op_net_x0;
  pilot <= logical1_y_net_x0;

  constant1: entity work.constant_1f05b15a2d
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_330e503d71
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_173d83e4a7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  constant4: entity work.constant_8207020ee3
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  logical1: entity work.logical_a6d07705dd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational4_op_net,
      d1(0) => relational5_op_net_x0,
      d2(0) => relational6_op_net,
      d3(0) => relational7_op_net,
      y(0) => logical1_y_net_x0
    );

  relational4: entity work.relational_931d61fb72
    port map (
      a => constant2_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational4_op_net
    );

  relational5: entity work.relational_931d61fb72
    port map (
      a => constant1_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational5_op_net_x0
    );

  relational6: entity work.relational_931d61fb72
    port map (
      a => constant4_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational6_op_net
    );

  relational7: entity work.relational_931d61fb72
    port map (
      a => constant3_op_net,
      b => subcarrier_index_op_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational7_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots/Pilot Gen/Scrambling LFSR"

entity scrambling_lfsr_entity_3984375e7e is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    q: out std_logic
  );
end scrambling_lfsr_entity_3984375e7e;

architecture structural of scrambling_lfsr_entity_3984375e7e is
  signal assert1_dout_net: std_logic;
  signal assert_dout_net: std_logic;
  signal ce_1_sg_x46: std_logic;
  signal clk_1_sg_x46: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x29: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register6_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x46 <= ce_1;
  clk_1_sg_x46 <= clk_1;
  logical1_y_net_x1 <= en;
  logical_y_net_x29 <= rst;
  q <= logical_y_net_x0;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register3_q_net,
      dout(0) => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register6_q_net,
      dout(0) => assert_dout_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      clr => '0',
      din(0) => logical_y_net_x29,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      clr => '0',
      din(0) => logical1_y_net_x1,
      en => "1",
      dout(0) => convert1_dout_net
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => assert_dout_net,
      d1(0) => assert1_dout_net,
      y(0) => logical_y_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register1_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register2_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register3_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register4_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => register5_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register6_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x46,
      clk => clk_1_sg_x46,
      d(0) => logical_y_net_x0,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots/Pilot Gen"

entity pilot_gen_entity_558a3ce157 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    reset: in std_logic; 
    sc_ind: in std_logic_vector(5 downto 0); 
    pilot_i: out std_logic_vector(11 downto 0); 
    pilot_valid: out std_logic
  );
end pilot_gen_entity_558a3ce157;

architecture structural of pilot_gen_entity_558a3ce157 is
  signal ce_1_sg_x47: std_logic;
  signal clk_1_sg_x47: std_logic;
  signal constant1_op_net: std_logic_vector(11 downto 0);
  signal constant5_op_net: std_logic_vector(11 downto 0);
  signal delay_q_net: std_logic_vector(5 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x30: std_logic;
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal relational1_op_net_x0: std_logic;
  signal relational5_op_net_x0: std_logic;
  signal subcarrier_index_op_net_x2: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x47 <= ce_1;
  clk_1_sg_x47 <= clk_1;
  logical_y_net_x30 <= reset;
  subcarrier_index_op_net_x2 <= sc_ind;
  pilot_i <= mux1_y_net_x0;
  pilot_valid <= logical1_y_net_x2;

  constant1: entity work.constant_e054d850c5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant5: entity work.constant_9127ce6619
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 6
    )
    port map (
      ce => ce_1_sg_x47,
      clk => clk_1_sg_x47,
      d => subcarrier_index_op_net_x2,
      en => '1',
      rst => '1',
      q => delay_q_net
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational5_op_net_x0,
      d1(0) => logical_y_net_x0,
      y(0) => logical_y_net
    );

  mux1: entity work.mux_4de2214a42
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant5_op_net,
      d1 => constant1_op_net,
      sel(0) => logical_y_net,
      y => mux1_y_net_x0
    );

  pilot_selection_93fec99adc: entity work.pilot_selection_entity_93fec99adc
    port map (
      sc_ind => subcarrier_index_op_net_x2,
      negate => relational5_op_net_x0,
      pilot => logical1_y_net_x2
    );

  posedge_ee6e94f233: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x47,
      clk_1 => clk_1_sg_x47,
      d => relational1_op_net_x0,
      q => logical1_y_net_x1
    );

  relational1: entity work.relational_47932db5b1
    port map (
      a => subcarrier_index_op_net_x2,
      b => delay_q_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  scrambling_lfsr_3984375e7e: entity work.scrambling_lfsr_entity_3984375e7e
    port map (
      ce_1 => ce_1_sg_x47,
      clk_1 => clk_1_sg_x47,
      en => logical1_y_net_x1,
      rst => logical_y_net_x30,
      q => logical_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots/Subcarrier Index Count"

entity subcarrier_index_count_entity_16356605e7 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    regtx_num_sc: in std_logic_vector(7 downto 0); 
    reset: in std_logic; 
    last: out std_logic; 
    sc_ind: out std_logic_vector(5 downto 0)
  );
end subcarrier_index_count_entity_16356605e7;

architecture structural of subcarrier_index_count_entity_16356605e7 is
  signal addsub_s_net: std_logic_vector(8 downto 0);
  signal b_7_0_y_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x52: std_logic;
  signal clk_1_sg_x52: std_logic;
  signal constant1_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net: std_logic;
  signal logical_y_net_x32: std_logic;
  signal relational3_op_net: std_logic;
  signal subcarrier_index_op_net_x3: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x52 <= ce_1;
  clk_1_sg_x52 <= clk_1;
  logical1_y_net_x1 <= en;
  b_7_0_y_net_x1 <= regtx_num_sc;
  logical_y_net_x32 <= reset;
  last <= logical1_y_net_x2;
  sc_ind <= subcarrier_index_op_net_x3;

  addsub: entity work.xladdsub_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 8,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 1,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 9,
      core_name0 => "addsb_11_0_a52ead9b8a3c1e76",
      extra_registers => 0,
      full_s_arith => 2,
      full_s_width => 9,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlSigned,
      s_bin_pt => 0,
      s_width => 9
    )
    port map (
      a => b_7_0_y_net_x1,
      b(0) => constant1_op_net,
      ce => ce_1_sg_x52,
      clk => clk_1_sg_x52,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => logical1_y_net_x1,
      y(0) => logical1_y_net_x2
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x32,
      d1(0) => logical1_y_net_x2,
      y(0) => logical2_y_net
    );

  relational3: entity work.relational_1834ac00b4
    port map (
      a => addsub_s_net,
      b => subcarrier_index_op_net_x3,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  subcarrier_index: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_f068fb73312ae1e5",
      op_arith => xlUnsigned,
      op_width => 6
    )
    port map (
      ce => ce_1_sg_x52,
      clk => clk_1_sg_x52,
      clr => '0',
      en(0) => logical1_y_net_x1,
      rst(0) => logical2_y_net,
      op => subcarrier_index_op_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/Control & Pilots"

entity \control___pilots_entity_f50034fe28\ is
  port (
    b_7_0: in std_logic_vector(7 downto 0); 
    bits_ready: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fifo_ready: in std_logic; 
    ppdu_tail_done: in std_logic; 
    tx_reset: in std_logic; 
    data: out std_logic; 
    data_sym_ind: out std_logic_vector(5 downto 0); 
    iq_sel: out std_logic_vector(1 downto 0); 
    iq_valid: out std_logic; 
    last_samp: out std_logic; 
    last_sym: out std_logic; 
    pilot_i: out std_logic_vector(11 downto 0)
  );
end \control___pilots_entity_f50034fe28\;

architecture structural of \control___pilots_entity_f50034fe28\ is
  signal axi_fifo_s_axis_tready_net_x1: std_logic;
  signal b_7_0_y_net_x2: std_logic_vector(7 downto 0);
  signal ce_1_sg_x53: std_logic;
  signal clk_1_sg_x53: std_logic;
  signal concat1_y_net: std_logic_vector(1 downto 0);
  signal delay1_q_net_x1: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x10: std_logic;
  signal delay3_q_net_x5: std_logic;
  signal delay3_q_net_x6: std_logic;
  signal delay4_q_net: std_logic;
  signal delay5_q_net_x0: std_logic_vector(1 downto 0);
  signal delay6_q_net_x0: std_logic_vector(11 downto 0);
  signal delay_q_net_x1: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical2_y_net: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x33: std_logic;
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal slice_y_net_x4: std_logic_vector(5 downto 0);
  signal subcarrier_index_op_net_x3: std_logic_vector(5 downto 0);

begin
  b_7_0_y_net_x2 <= b_7_0;
  delay2_q_net_x10 <= bits_ready;
  ce_1_sg_x53 <= ce_1;
  clk_1_sg_x53 <= clk_1;
  axi_fifo_s_axis_tready_net_x1 <= fifo_ready;
  delay3_q_net_x5 <= ppdu_tail_done;
  logical_y_net_x33 <= tx_reset;
  data <= delay2_q_net_x0;
  data_sym_ind <= slice_y_net_x4;
  iq_sel <= delay5_q_net_x0;
  iq_valid <= delay_q_net_x1;
  last_samp <= delay1_q_net_x1;
  last_sym <= delay3_q_net_x6;
  pilot_i <= delay6_q_net_x0;

  concat1: entity work.concat_32afb77cd2
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => relational1_op_net_x0,
      in1(0) => logical1_y_net_x2,
      y => concat1_y_net
    );

  data_sc_map_0f52ca1546: entity work.data_sc_map_entity_0f52ca1546
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      sc_ind => subcarrier_index_op_net_x3,
      data_sym_ind => slice_y_net_x4,
      data_sym_valid => relational1_op_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x1
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d(0) => logical1_y_net_x5,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x1
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d(0) => register2_q_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  delay3: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d(0) => logical2_y_net,
      en => '1',
      rst => '1',
      q(0) => delay3_q_net_x6
    );

  delay4: entity work.delay_0341f7be44
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d(0) => delay3_q_net_x5,
      q(0) => delay4_q_net
    );

  delay5: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 2
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d => concat1_y_net,
      en => '1',
      rst => '1',
      q => delay5_q_net_x0
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 12
    )
    port map (
      ce => ce_1_sg_x53,
      clk => clk_1_sg_x53,
      d => mux1_y_net_x0,
      en => '1',
      rst => '1',
      q => delay6_q_net_x0
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x33,
      d1(0) => logical1_y_net_x5,
      y(0) => logical_y_net_x0
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => axi_fifo_s_axis_tready_net_x1,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x5,
      d1(0) => delay4_q_net,
      y(0) => logical2_y_net
    );

  pilot_gen_558a3ce157: entity work.pilot_gen_entity_558a3ce157
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      reset => logical_y_net_x33,
      sc_ind => subcarrier_index_op_net_x3,
      pilot_i => mux1_y_net_x0,
      pilot_valid => logical1_y_net_x2
    );

  posedge1_45ac091708: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      d => logical_y_net_x0,
      q => logical1_y_net_x4
    );

  posedge_e39e2937a0: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      d => delay2_q_net_x10,
      q => logical1_y_net_x3
    );

  s_r_latch1_9fcc1a0be5: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      r => logical1_y_net_x4,
      s => logical1_y_net_x3,
      q => register2_q_net_x0
    );

  s_r_latch2_a5fc701055: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      r => logical_y_net_x33,
      s => logical1_y_net_x5,
      q => register2_q_net_x1
    );

  subcarrier_index_count_16356605e7: entity work.subcarrier_index_count_entity_16356605e7
    port map (
      ce_1 => ce_1_sg_x53,
      clk_1 => clk_1_sg_x53,
      en => logical1_y_net_x1,
      regtx_num_sc => b_7_0_y_net_x2,
      reset => logical_y_net_x33,
      last => logical1_y_net_x5,
      sc_ind => subcarrier_index_op_net_x3
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/QPSK/QPSK Int Addr"

entity qpsk_int_addr_entity_dd03169980 is
  port (
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    new_sym: in std_logic; 
    tx_reset: in std_logic; 
    wr_addr: out std_logic_vector(6 downto 0); 
    wr_offset: out std_logic
  );
end qpsk_int_addr_entity_dd03169980;

architecture structural of qpsk_int_addr_entity_dd03169980 is
  signal ce_1_sg_x56: std_logic;
  signal clk_1_sg_x56: std_logic;
  signal constant2_op_net: std_logic_vector(6 downto 0);
  signal counter_op_net: std_logic_vector(6 downto 0);
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x11: std_logic;
  signal delay_q_net_x7: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x35: std_logic;
  signal qpsk_int1_data_net_x0: std_logic_vector(6 downto 0);
  signal register2_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;

begin
  delay_q_net_x7 <= bit_valid;
  ce_1_sg_x56 <= ce_1;
  clk_1_sg_x56 <= clk_1;
  delay2_q_net_x11 <= new_sym;
  logical_y_net_x35 <= tx_reset;
  wr_addr <= qpsk_int1_data_net_x0;
  wr_offset <= delay2_q_net_x0;

  constant2: entity work.constant_011ca80190
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  counter: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 95,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_d24951bef2f0cdc9",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 7
    )
    port map (
      ce => ce_1_sg_x56,
      clk => clk_1_sg_x56,
      clr => '0',
      en(0) => delay_q_net_x7,
      rst(0) => logical1_y_net,
      op => counter_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x56,
      clk => clk_1_sg_x56,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  logical1: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x35,
      d1(0) => delay2_q_net_x11,
      d2(0) => logical1_y_net_x1,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x7,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  osc_0375f0cbbe: entity work.osc_entity_4b2508a4db
    port map (
      ce_1 => ce_1_sg_x56,
      clk_1 => clk_1_sg_x56,
      en => logical1_y_net_x1,
      r => logical_y_net_x35,
      q => register2_q_net_x0
    );

  posedge_7727a40979: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x56,
      clk_1 => clk_1_sg_x56,
      d => logical2_y_net_x0,
      q => logical1_y_net_x1
    );

  qpsk_int1: entity work.xlsprom_wlan_phy_tx_pmd
    generic map (
      c_address_width => 7,
      c_width => 7,
      core_name0 => "bmg_72_3628803596b5ca22",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x56,
      clk => clk_1_sg_x56,
      en => "1",
      rst => "0",
      data => qpsk_int1_data_net_x0
    );

  relational2: entity work.relational_9a3978c602
    port map (
      a => counter_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/QPSK"

entity qpsk_entity_07b9523b2d is
  port (
    bit_tdata: in std_logic; 
    bit_tvalid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_sym_addr: in std_logic_vector(5 downto 0); 
    logical: in std_logic; 
    new_sym: in std_logic; 
    x2b_data: out std_logic_vector(1 downto 0)
  );
end qpsk_entity_07b9523b2d;

architecture structural of qpsk_entity_07b9523b2d is
  signal bit_memory1_doutb_net_x0: std_logic_vector(1 downto 0);
  signal ce_1_sg_x57: std_logic;
  signal clk_1_sg_x57: std_logic;
  signal concat1_y_net: std_logic_vector(7 downto 0);
  signal concat2_y_net: std_logic_vector(6 downto 0);
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic;
  signal delay2_q_net: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x12: std_logic;
  signal delay6_q_net: std_logic;
  signal delay_q_net_x8: std_logic;
  signal inverter_op_net: std_logic;
  signal logical_y_net_x36: std_logic;
  signal mux_y_net_x3: std_logic;
  signal qpsk_int1_data_net_x0: std_logic_vector(6 downto 0);
  signal slice_y_net_x5: std_logic_vector(5 downto 0);

begin
  mux_y_net_x3 <= bit_tdata;
  delay_q_net_x8 <= bit_tvalid;
  ce_1_sg_x57 <= ce_1;
  clk_1_sg_x57 <= clk_1;
  slice_y_net_x5 <= data_sym_addr;
  logical_y_net_x36 <= logical;
  delay2_q_net_x12 <= new_sym;
  x2b_data <= bit_memory1_doutb_net_x0;

  bit_memory1: entity work.xldpram_wlan_phy_tx_pmd
    generic map (
      c_address_width_a => 8,
      c_address_width_b => 7,
      c_width_a => 1,
      c_width_b => 2,
      core_name0 => "bmg_72_376dc060ca4075f2",
      latency => 1
    )
    port map (
      a_ce => ce_1_sg_x57,
      a_clk => clk_1_sg_x57,
      addra => concat1_y_net,
      addrb => concat2_y_net,
      b_ce => ce_1_sg_x57,
      b_clk => clk_1_sg_x57,
      dina(0) => delay6_q_net,
      dinb => constant1_op_net,
      ena => "1",
      enb => "1",
      rsta => "0",
      rstb => "0",
      wea(0) => delay2_q_net,
      web(0) => constant2_op_net,
      doutb => bit_memory1_doutb_net_x0
    );

  concat1: entity work.concat_83e473517e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => delay2_q_net_x0,
      in1 => qpsk_int1_data_net_x0,
      y => concat1_y_net
    );

  concat2: entity work.concat_c6a9b6687e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => inverter_op_net,
      in1 => slice_y_net_x5,
      y => concat2_y_net
    );

  constant1: entity work.constant_cda50df78a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  delay2: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => delay_q_net_x8,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net
    );

  delay6: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      d(0) => mux_y_net_x3,
      en => '1',
      rst => '1',
      q(0) => delay6_q_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x57,
      clk => clk_1_sg_x57,
      clr => '0',
      ip(0) => delay2_q_net_x0,
      op(0) => inverter_op_net
    );

  qpsk_int_addr_dd03169980: entity work.qpsk_int_addr_entity_dd03169980
    port map (
      bit_valid => delay_q_net_x8,
      ce_1 => ce_1_sg_x57,
      clk_1 => clk_1_sg_x57,
      new_sym => delay2_q_net_x12,
      tx_reset => logical_y_net_x36,
      wr_addr => qpsk_int1_data_net_x0,
      wr_offset => delay2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate/QPSK Mod"

entity qpsk_mod_entity_eb137744eb is
  port (
    b_1_0: in std_logic_vector(1 downto 0); 
    i: out std_logic_vector(11 downto 0); 
    q: out std_logic_vector(11 downto 0)
  );
end qpsk_mod_entity_eb137744eb;

architecture structural of qpsk_mod_entity_eb137744eb is
  signal bit_memory1_doutb_net_x1: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(11 downto 0);
  signal constant3_op_net: std_logic_vector(11 downto 0);
  signal lsb_1_y_net: std_logic;
  signal lsb_y_net: std_logic;
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);

begin
  bit_memory1_doutb_net_x1 <= b_1_0;
  i <= mux_y_net_x0;
  q <= mux1_y_net_x0;

  constant2: entity work.constant_2a9931b0e7
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant3: entity work.constant_40d4599892
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => bit_memory1_doutb_net_x1,
      y(0) => lsb_y_net
    );

  lsb_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 2,
      y_width => 1
    )
    port map (
      x => bit_memory1_doutb_net_x1,
      y(0) => lsb_1_y_net
    );

  mux: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => lsb_y_net,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_c3e1ddb86e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant2_op_net,
      d1 => constant3_op_net,
      sel(0) => lsb_1_y_net,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Interleave & Modulate"

entity \interleave___modulate_entity_1e78258d30\ is
  port (
    b_7_0: in std_logic_vector(7 downto 0); 
    bit: in std_logic; 
    bit_source: in std_logic; 
    bit_source_x0: in std_logic_vector(8 downto 0); 
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fifo_in_ready: in std_logic; 
    logical: in std_logic; 
    signal_mod_sel: in std_logic_vector(1 downto 0); 
    last_sym: out std_logic; 
    x_i: out std_logic_vector(11 downto 0); 
    x_iq_last: out std_logic; 
    x_iq_valid: out std_logic; 
    x_q: out std_logic_vector(11 downto 0)
  );
end \interleave___modulate_entity_1e78258d30\;

architecture structural of \interleave___modulate_entity_1e78258d30\ is
  signal axi_fifo_s_axis_tready_net_x2: std_logic;
  signal b_2_1_y_net_x1: std_logic_vector(1 downto 0);
  signal b_7_0_y_net_x3: std_logic_vector(7 downto 0);
  signal bit_memory1_doutb_net_x1: std_logic_vector(3 downto 0);
  signal bit_memory1_doutb_net_x2: std_logic_vector(1 downto 0);
  signal bit_memory_doutb_net_x1: std_logic;
  signal ce_1_sg_x58: std_logic;
  signal clk_1_sg_x58: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal constant4_op_net_x0: std_logic_vector(11 downto 0);
  signal constant5_op_net: std_logic_vector(11 downto 0);
  signal constant6_op_net: std_logic_vector(11 downto 0);
  signal convert2_dout_net: std_logic;
  signal convert2_dout_net_x5: std_logic_vector(8 downto 0);
  signal delay1_q_net_x2: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal delay2_q_net_x12: std_logic;
  signal delay3_q_net_x7: std_logic;
  signal delay3_q_net_x8: std_logic;
  signal delay5_q_net_x0: std_logic_vector(1 downto 0);
  signal delay6_q_net_x0: std_logic_vector(11 downto 0);
  signal delay_q_net_x10: std_logic;
  signal delay_q_net_x9: std_logic;
  signal logical2_y_net: std_logic_vector(1 downto 0);
  signal logical_y_net_x37: std_logic;
  signal mux1_y_net: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(11 downto 0);
  signal mux1_y_net_x1: std_logic_vector(11 downto 0);
  signal mux1_y_net_x2: std_logic_vector(11 downto 0);
  signal mux2_y_net: std_logic_vector(11 downto 0);
  signal mux3_y_net_x1: std_logic_vector(11 downto 0);
  signal mux4_y_net_x1: std_logic_vector(11 downto 0);
  signal mux_y_net_x0: std_logic_vector(11 downto 0);
  signal mux_y_net_x1: std_logic_vector(11 downto 0);
  signal mux_y_net_x2: std_logic_vector(11 downto 0);
  signal mux_y_net_x3: std_logic_vector(11 downto 0);
  signal mux_y_net_x5: std_logic;
  signal slice_y_net_x3: std_logic_vector(5 downto 0);
  signal slice_y_net_x5: std_logic_vector(5 downto 0);

begin
  b_7_0_y_net_x3 <= b_7_0;
  mux_y_net_x5 <= bit;
  delay3_q_net_x7 <= bit_source;
  convert2_dout_net_x5 <= bit_source_x0;
  delay_q_net_x9 <= bit_valid;
  ce_1_sg_x58 <= ce_1;
  clk_1_sg_x58 <= clk_1;
  axi_fifo_s_axis_tready_net_x2 <= fifo_in_ready;
  logical_y_net_x37 <= logical;
  b_2_1_y_net_x1 <= signal_mod_sel;
  last_sym <= delay3_q_net_x8;
  x_i <= mux3_y_net_x1;
  x_iq_last <= delay1_q_net_x2;
  x_iq_valid <= delay_q_net_x10;
  x_q <= mux4_y_net_x1;

  bpsk_ba0b27afd0: entity work.bpsk_entity_ba0b27afd0
    port map (
      bit_tdata => mux_y_net_x5,
      bit_tvalid => delay_q_net_x9,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      data_sym_addr => slice_y_net_x5,
      logical => logical_y_net_x37,
      new_sym => delay2_q_net_x12,
      x1b_data => bit_memory_doutb_net_x1
    );

  bpsk_mod_9dd399b8d9: entity work.bpsk_mod_entity_9dd399b8d9
    port map (
      b_0 => bit_memory_doutb_net_x1,
      i => mux_y_net_x2,
      q => constant4_op_net_x0
    );

  coded_bit_counter_bb3901367b: entity work.coded_bit_counter_entity_bb3901367b
    port map (
      bit_valid => delay_q_net_x9,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      data_n_cbps => convert2_dout_net_x5,
      tx_reset => logical_y_net_x37,
      bits_ready => delay2_q_net_x12
    );

  concat: entity work.concat_e6f5ee726b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => convert2_dout_net,
      in1(0) => convert2_dout_net,
      y => concat_y_net
    );

  constant5: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant5_op_net
    );

  constant6: entity work.constant_fd28b32bf8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant6_op_net
    );

  control_pilots_f50034fe28: entity work.\control___pilots_entity_f50034fe28\
    port map (
      b_7_0 => b_7_0_y_net_x3,
      bits_ready => delay2_q_net_x12,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      fifo_ready => axi_fifo_s_axis_tready_net_x2,
      ppdu_tail_done => delay3_q_net_x7,
      tx_reset => logical_y_net_x37,
      data => delay2_q_net_x0,
      data_sym_ind => slice_y_net_x5,
      iq_sel => delay5_q_net_x0,
      iq_valid => delay_q_net_x10,
      last_samp => delay1_q_net_x2,
      last_sym => delay3_q_net_x8,
      pilot_i => delay6_q_net_x0
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x58,
      clk => clk_1_sg_x58,
      clr => '0',
      din(0) => delay2_q_net_x0,
      en => "1",
      dout(0) => convert2_dout_net
    );

  logical2: entity work.logical_33c9a0c803
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => b_2_1_y_net_x1,
      d1 => concat_y_net,
      y => logical2_y_net
    );

  mux1: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => mux_y_net_x2,
      d1 => mux_y_net_x3,
      d2 => mux_y_net_x0,
      d3 => mux_y_net_x1,
      sel => logical2_y_net,
      y => mux1_y_net
    );

  mux2: entity work.mux_192c5da026
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant4_op_net_x0,
      d1 => mux1_y_net_x2,
      d2 => mux1_y_net_x0,
      d3 => mux1_y_net_x1,
      sel => logical2_y_net,
      y => mux2_y_net
    );

  mux3: entity work.mux_e5a9964709
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant6_op_net,
      d1 => delay6_q_net_x0,
      d2 => mux1_y_net,
      sel => delay5_q_net_x0,
      y => mux3_y_net_x1
    );

  mux4: entity work.mux_e5a9964709
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => constant5_op_net,
      d1 => constant5_op_net,
      d2 => mux2_y_net,
      sel => delay5_q_net_x0,
      y => mux4_y_net_x1
    );

  qpsk_07b9523b2d: entity work.qpsk_entity_07b9523b2d
    port map (
      bit_tdata => mux_y_net_x5,
      bit_tvalid => delay_q_net_x9,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      data_sym_addr => slice_y_net_x5,
      logical => logical_y_net_x37,
      new_sym => delay2_q_net_x12,
      x2b_data => bit_memory1_doutb_net_x2
    );

  qpsk_mod_eb137744eb: entity work.qpsk_mod_entity_eb137744eb
    port map (
      b_1_0 => bit_memory1_doutb_net_x2,
      i => mux_y_net_x3,
      q => mux1_y_net_x2
    );

  x16_qam_381a479990: entity work.x16_qam_entity_381a479990
    port map (
      bit_tdata => mux_y_net_x5,
      bit_tvalid => delay_q_net_x9,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      data_sym_addr => slice_y_net_x5,
      logical => logical_y_net_x37,
      new_sym => delay2_q_net_x12,
      x4b_data => bit_memory1_doutb_net_x1
    );

  x16qam_mod_cce570a88c: entity work.x16qam_mod_entity_cce570a88c
    port map (
      b_3_0 => bit_memory1_doutb_net_x1,
      i => mux_y_net_x0,
      q => mux1_y_net_x0
    );

  x64_qam_35dea913c2: entity work.x64_qam_entity_35dea913c2
    port map (
      bit_tdata => mux_y_net_x5,
      bit_tvalid => delay_q_net_x9,
      ce_1 => ce_1_sg_x58,
      clk_1 => clk_1_sg_x58,
      data_sym_addr => slice_y_net_x5,
      logical => logical_y_net_x37,
      new_sym => delay2_q_net_x12,
      x6b_data => slice_y_net_x3
    );

  x64qam_mod_e734ca01a6: entity work.x64qam_mod_entity_e734ca01a6
    port map (
      b_5_0 => slice_y_net_x3,
      i => mux_y_net_x1,
      q => mux1_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/DAC Outputs"

entity dac_outputs_entity_fec48642b9 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    i: in std_logic_vector(11 downto 0); 
    q: in std_logic_vector(11 downto 0); 
    regtx_anta_tx_en: in std_logic; 
    regtx_antb_tx_en: in std_logic; 
    register1_x0: out std_logic_vector(11 downto 0); 
    register2_x0: out std_logic_vector(11 downto 0); 
    register3_x0: out std_logic_vector(11 downto 0); 
    register_x1: out std_logic_vector(11 downto 0)
  );
end dac_outputs_entity_fec48642b9;

architecture structural of dac_outputs_entity_fec48642b9 is
  signal b_2_y_net: std_logic;
  signal b_3_y_net: std_logic;
  signal ce_1_sg_x59: std_logic;
  signal clk_1_sg_x59: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical_y_net: std_logic;
  signal mult1_p_net_x0: std_logic_vector(11 downto 0);
  signal mult_p_net_x0: std_logic_vector(11 downto 0);
  signal register1_q_net_x0: std_logic_vector(11 downto 0);
  signal register2_q_net_x0: std_logic_vector(11 downto 0);
  signal register3_q_net_x0: std_logic_vector(11 downto 0);
  signal register_q_net_x0: std_logic_vector(11 downto 0);

begin
  ce_1_sg_x59 <= ce_1;
  clk_1_sg_x59 <= clk_1;
  logical1_y_net_x1 <= en;
  mult_p_net_x0 <= i;
  mult1_p_net_x0 <= q;
  b_2_y_net <= regtx_anta_tx_en;
  b_3_y_net <= regtx_antb_tx_en;
  register1_x0 <= register1_q_net_x0;
  register2_x0 <= register2_q_net_x0;
  register3_x0 <= register3_q_net_x0;
  register_x1 <= register_q_net_x0;

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      ip(0) => logical_y_net,
      op(0) => inverter1_op_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      clr => '0',
      ip(0) => logical1_y_net,
      op(0) => inverter2_op_net
    );

  logical: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => b_2_y_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => b_3_y_net,
      y(0) => logical1_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      d => mult1_p_net_x0,
      en => "1",
      rst(0) => inverter1_op_net,
      q => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      d => mult_p_net_x0,
      en => "1",
      rst(0) => inverter2_op_net,
      q => register2_q_net_x0
    );

  register3: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      d => mult1_p_net_x0,
      en => "1",
      rst(0) => inverter2_op_net,
      q => register3_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x59,
      clk => clk_1_sg_x59,
      d => mult_p_net_x0,
      en => "1",
      rst(0) => inverter1_op_net,
      q => register_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/FIFO/I/Q Concat"

entity q_concat_entity_9872452a0b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    q: in std_logic_vector(15 downto 0); 
    iq: out std_logic_vector(31 downto 0)
  );
end q_concat_entity_9872452a0b;

architecture structural of q_concat_entity_9872452a0b is
  signal ce_1_sg_x60: std_logic;
  signal clk_1_sg_x60: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert1_dout_net: std_logic_vector(15 downto 0);
  signal convert_dout_net: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x60 <= ce_1;
  clk_1_sg_x60 <= clk_1;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2 <= i;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2 <= q;
  iq <= concat_y_net_x0;

  concat: entity work.concat_a369e00c6b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => reinterpret_output_port_net,
      in1 => reinterpret1_output_port_net,
      y => concat_y_net_x0
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      din => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x2,
      en => "1",
      dout => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 2,
      din_bin_pt => 15,
      din_width => 16,
      dout_arith => 2,
      dout_bin_pt => 15,
      dout_width => 16,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x60,
      clk => clk_1_sg_x60,
      clr => '0',
      din => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x2,
      en => "1",
      dout => convert1_dout_net
    );

  reinterpret: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert_dout_net,
      output_port => reinterpret_output_port_net
    );

  reinterpret1: entity work.reinterpret_7025463ea8
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => convert1_dout_net,
      output_port => reinterpret1_output_port_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/FIFO"

entity fifo_entity_ed2bc31ace is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_i: in std_logic_vector(15 downto 0); 
    fft_q: in std_logic_vector(15 downto 0); 
    rd: in std_logic; 
    reset: in std_logic; 
    tx_reset: in std_logic; 
    write: in std_logic; 
    i: out std_logic_vector(15 downto 0); 
    occ: out std_logic_vector(7 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end fifo_entity_ed2bc31ace;

architecture structural of fifo_entity_ed2bc31ace is
  signal ce_1_sg_x61: std_logic;
  signal clk_1_sg_x61: std_logic;
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal convert2_dout_net: std_logic;
  signal delay1_q_net: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x3: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x3: std_logic_vector(15 downto 0);
  signal fifo_dcount_net_x2: std_logic_vector(7 downto 0);
  signal fifo_dout_net_x0: std_logic_vector(31 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical4_y_net: std_logic;
  signal logical4_y_net_x1: std_logic;
  signal logical_y_net_x38: std_logic;
  signal reinterpret2_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x61 <= ce_1;
  clk_1_sg_x61 <= clk_1;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x3 <= fft_i;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x3 <= fft_q;
  logical2_y_net_x0 <= rd;
  logical1_y_net_x0 <= reset;
  logical_y_net_x38 <= tx_reset;
  logical4_y_net_x1 <= write;
  i <= reinterpret2_output_port_net_x1;
  occ <= fifo_dcount_net_x2;
  q <= reinterpret3_output_port_net_x1;

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      clr => '0',
      din(0) => logical1_y_net_x0,
      en => "1",
      dout(0) => convert2_dout_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 12,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      d(0) => logical_y_net_x38,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  fifo: entity work.xlfifogen_wlan_phy_tx_pmd
    generic map (
      core_name0 => "fifo_fg92_6a1156e8dc43a711",
      data_count_width => 8,
      data_width => 32,
      has_ae => 0,
      has_af => 0,
      percent_full_width => 1
    )
    port map (
      ce => ce_1_sg_x61,
      clk => clk_1_sg_x61,
      din => concat_y_net_x0,
      en => '1',
      re => logical2_y_net_x0,
      re_ce => ce_1_sg_x61,
      rst => logical4_y_net,
      we => logical4_y_net_x1,
      we_ce => ce_1_sg_x61,
      dcount => fifo_dcount_net_x2,
      dout => fifo_dout_net_x0
    );

  logical4: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay1_q_net,
      d1(0) => convert2_dout_net,
      y(0) => logical4_y_net
    );

  q_concat_9872452a0b: entity work.q_concat_entity_9872452a0b
    port map (
      ce_1 => ce_1_sg_x61,
      clk_1 => clk_1_sg_x61,
      i => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x3,
      q => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x3,
      iq => concat_y_net_x0
    );

  q_slice_a49b8b75e5: entity work.q_slice_entity_10657a6c34
    port map (
      iq => fifo_dout_net_x0,
      i => reinterpret2_output_port_net_x1,
      q => reinterpret3_output_port_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/Preamble Gen"

entity preamble_gen_entity_c25e867a97 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    rd_en: in std_logic; 
    tx_reset: in std_logic; 
    tx_running: in std_logic; 
    done: out std_logic; 
    early_done: out std_logic; 
    i: out std_logic_vector(15 downto 0); 
    q: out std_logic_vector(15 downto 0)
  );
end preamble_gen_entity_c25e867a97;

architecture structural of preamble_gen_entity_c25e867a97 is
  signal ce_1_sg_x63: std_logic;
  signal clk_1_sg_x63: std_logic;
  signal constant3_op_net: std_logic_vector(8 downto 0);
  signal convert2_dout_net_x3: std_logic;
  signal counter_op_net: std_logic_vector(8 downto 0);
  signal delay4_q_net: std_logic;
  signal inverter1_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical_y_net_x39: std_logic;
  signal preamble_i_data_net: std_logic_vector(15 downto 0);
  signal preamble_q_data_net: std_logic_vector(15 downto 0);
  signal register1_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x2: std_logic_vector(15 downto 0);
  signal register3_q_net_x0: std_logic_vector(15 downto 0);
  signal register_q_net_x0: std_logic;
  signal relational2_op_net: std_logic;

begin
  ce_1_sg_x63 <= ce_1;
  clk_1_sg_x63 <= clk_1;
  convert2_dout_net_x3 <= rd_en;
  logical_y_net_x39 <= tx_reset;
  register2_q_net_x1 <= tx_running;
  done <= register1_q_net_x0;
  early_done <= register_q_net_x0;
  i <= register2_q_net_x2;
  q <= register3_q_net_x0;

  constant3: entity work.constant_0512fd5e4c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  counter: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_36e2bb554c95560d",
      op_arith => xlUnsigned,
      op_width => 9
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => delay4_q_net,
      op => counter_op_net
    );

  delay4: entity work.xldelay
    generic map (
      latency => 4,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d(0) => logical_y_net_x39,
      en => '1',
      rst => '1',
      q(0) => delay4_q_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      clr => '0',
      ip(0) => relational2_op_net,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x1,
      d1(0) => convert2_dout_net_x3,
      d2(0) => relational2_op_net,
      y(0) => logical1_y_net
    );

  preamble_i: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 9,
      c_address_width => 9,
      c_width => 16,
      core_name0 => "dmg_72_28ec6cac12d9767d",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      en => "1",
      data => preamble_i_data_net
    );

  preamble_q: entity work.xlsprom_dist_wlan_phy_tx_pmd
    generic map (
      addr_width => 9,
      c_address_width => 9,
      c_width => 16,
      core_name0 => "dmg_72_140171b6b191950b",
      latency => 1
    )
    port map (
      addr => counter_op_net,
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      en => "1",
      data => preamble_q_data_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d(0) => register_q_net_x0,
      en(0) => convert2_dout_net_x3,
      rst(0) => delay4_q_net,
      q(0) => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d => preamble_i_data_net,
      en(0) => convert2_dout_net_x3,
      rst(0) => delay4_q_net,
      q => register2_q_net_x2
    );

  register3: entity work.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d => preamble_q_data_net,
      en(0) => convert2_dout_net_x3,
      rst(0) => delay4_q_net,
      q => register3_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x63,
      clk => clk_1_sg_x63,
      d(0) => inverter1_op_net,
      en(0) => convert2_dout_net_x3,
      rst(0) => delay4_q_net,
      q(0) => register_q_net_x0
    );

  relational2: entity work.relational_82fb466a8b
    port map (
      a => counter_op_net,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs/Scaling"

entity scaling_entity_a269710a35 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    i: in std_logic_vector(15 downto 0); 
    preamble: in std_logic; 
    q: in std_logic_vector(15 downto 0); 
    regtx_scaling_payload: in std_logic_vector(15 downto 0); 
    regtx_scaling_preamble: in std_logic_vector(15 downto 0); 
    i_x0: out std_logic_vector(11 downto 0); 
    q_x0: out std_logic_vector(11 downto 0)
  );
end scaling_entity_a269710a35;

architecture structural of scaling_entity_a269710a35 is
  signal ce_1_sg_x66: std_logic;
  signal clk_1_sg_x66: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal mult1_p_net_x1: std_logic_vector(11 downto 0);
  signal mult_p_net_x1: std_logic_vector(11 downto 0);
  signal mux1_y_net_x0: std_logic_vector(15 downto 0);
  signal mux1_y_net_x1: std_logic_vector(15 downto 0);
  signal mux_y_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret1_output_port_net_x0: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net_x0: std_logic_vector(15 downto 0);

begin
  ce_1_sg_x66 <= ce_1;
  clk_1_sg_x66 <= clk_1;
  mux_y_net_x0 <= i;
  delay1_q_net_x0 <= preamble;
  mux1_y_net_x1 <= q;
  reinterpret1_output_port_net_x0 <= regtx_scaling_payload;
  reinterpret_output_port_net_x0 <= regtx_scaling_preamble;
  i_x0 <= mult_p_net_x1;
  q_x0 <= mult1_p_net_x1;

  mult: entity work.xlmult_wlan_phy_tx_pmd
    generic map (
      a_arith => xlSigned,
      a_bin_pt => 15,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 12,
      b_width => 16,
      c_a_type => 0,
      c_a_width => 16,
      c_b_type => 1,
      c_b_width => 16,
      c_baat => 16,
      c_output_width => 32,
      c_type => 0,
      core_name0 => "mult_11_2_f2bb5a57782af7d9",
      extra_registers => 1,
      multsign => 2,
      overflow => 2,
      p_arith => xlSigned,
      p_bin_pt => 11,
      p_width => 12,
      quantization => 1
    )
    port map (
      a => mux_y_net_x0,
      b => mux1_y_net_x0,
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      clr => '0',
      core_ce => ce_1_sg_x66,
      core_clk => clk_1_sg_x66,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult_p_net_x1
    );

  mult1: entity work.xlmult_wlan_phy_tx_pmd
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 12,
      a_width => 16,
      b_arith => xlSigned,
      b_bin_pt => 15,
      b_width => 16,
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 0,
      c_b_width => 16,
      c_baat => 16,
      c_output_width => 32,
      c_type => 0,
      core_name0 => "mult_11_2_414c0fa5acc33f35",
      extra_registers => 1,
      multsign => 2,
      overflow => 2,
      p_arith => xlSigned,
      p_bin_pt => 11,
      p_width => 12,
      quantization => 1
    )
    port map (
      a => mux1_y_net_x0,
      b => mux1_y_net_x1,
      ce => ce_1_sg_x66,
      clk => clk_1_sg_x66,
      clr => '0',
      core_ce => ce_1_sg_x66,
      core_clk => clk_1_sg_x66,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult1_p_net_x1
    );

  mux1: entity work.mux_a54904b290
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => reinterpret1_output_port_net_x0,
      d1 => reinterpret_output_port_net_x0,
      sel(0) => delay1_q_net_x0,
      y => mux1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Preamble & Outputs"

entity \preamble___outputs_entity_82fcc722dc\ is
  port (
    b_2: in std_logic; 
    b_3: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    fft_i: in std_logic_vector(15 downto 0); 
    fft_i_q_valid: in std_logic; 
    fft_q: in std_logic_vector(15 downto 0); 
    last_sym: in std_logic; 
    reinterpret: in std_logic_vector(15 downto 0); 
    reinterpret1: in std_logic_vector(15 downto 0); 
    tx_iq_samp_ce: in std_logic; 
    tx_reset: in std_logic; 
    tx_start: in std_logic; 
    dac_outputs: out std_logic_vector(11 downto 0); 
    dac_outputs_x0: out std_logic_vector(11 downto 0); 
    dac_outputs_x1: out std_logic_vector(11 downto 0); 
    dac_outputs_x2: out std_logic_vector(11 downto 0); 
    last_samp_output_to_dacs: out std_logic; 
    output_fifo_occ: out std_logic_vector(7 downto 0)
  );
end \preamble___outputs_entity_82fcc722dc\;

architecture structural of \preamble___outputs_entity_82fcc722dc\ is
  signal b_2_y_net_x0: std_logic;
  signal b_3_y_net_x0: std_logic;
  signal ce_1_sg_x67: std_logic;
  signal clk_1_sg_x67: std_logic;
  signal constant2_op_net: std_logic;
  signal convert2_dout_net_x4: std_logic;
  signal delay1_q_net_x0: std_logic;
  signal delay2_q_net_x0: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2: std_logic;
  signal fifo_dcount_net_x3: std_logic_vector(7 downto 0);
  signal inverter1_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net_x1: std_logic;
  signal logical_y_net_x3: std_logic;
  signal logical_y_net_x4: std_logic;
  signal logical_y_net_x42: std_logic;
  signal mult1_p_net_x1: std_logic_vector(11 downto 0);
  signal mult_p_net_x1: std_logic_vector(11 downto 0);
  signal mux1_y_net_x1: std_logic_vector(15 downto 0);
  signal mux_y_net_x0: std_logic_vector(15 downto 0);
  signal register1_q_net_x1: std_logic;
  signal register1_q_net_x2: std_logic_vector(11 downto 0);
  signal register2_q_net_x2: std_logic_vector(15 downto 0);
  signal register2_q_net_x3: std_logic;
  signal register2_q_net_x4: std_logic;
  signal register2_q_net_x5: std_logic_vector(11 downto 0);
  signal register3_q_net_x1: std_logic_vector(15 downto 0);
  signal register3_q_net_x2: std_logic_vector(11 downto 0);
  signal register_q_net_x1: std_logic;
  signal register_q_net_x2: std_logic_vector(11 downto 0);
  signal reinterpret1_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x1: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net_x1: std_logic_vector(15 downto 0);
  signal relational1_op_net: std_logic;

begin
  b_2_y_net_x0 <= b_2;
  b_3_y_net_x0 <= b_3;
  ce_1_sg_x67 <= ce_1;
  clk_1_sg_x67 <= clk_1;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4 <= fft_i;
  fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2 <= fft_i_q_valid;
  fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4 <= fft_q;
  logical_y_net_x3 <= last_sym;
  reinterpret_output_port_net_x1 <= reinterpret;
  reinterpret1_output_port_net_x1 <= reinterpret1;
  convert2_dout_net_x4 <= tx_iq_samp_ce;
  logical_y_net_x42 <= tx_reset;
  logical_y_net_x4 <= tx_start;
  dac_outputs <= register_q_net_x2;
  dac_outputs_x0 <= register1_q_net_x2;
  dac_outputs_x1 <= register2_q_net_x5;
  dac_outputs_x2 <= register3_q_net_x2;
  last_samp_output_to_dacs <= delay2_q_net_x0;
  output_fifo_occ <= fifo_dcount_net_x3;

  constant2: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant2_op_net
    );

  dac_outputs_fec48642b9: entity work.dac_outputs_entity_fec48642b9
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      en => logical1_y_net_x1,
      i => mult_p_net_x1,
      q => mult1_p_net_x1,
      regtx_anta_tx_en => b_2_y_net_x0,
      regtx_antb_tx_en => b_3_y_net_x0,
      register1_x0 => register1_q_net_x2,
      register2_x0 => register2_q_net_x5,
      register3_x0 => register3_q_net_x2,
      register_x1 => register_q_net_x2
    );

  delay1: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      d(0) => register1_q_net_x1,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net_x0
    );

  delay2: entity work.xldelay
    generic map (
      latency => 12,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      d(0) => logical3_y_net,
      en => '1',
      rst => '1',
      q(0) => delay2_q_net_x0
    );

  fifo_ed2bc31ace: entity work.fifo_entity_ed2bc31ace
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      fft_i => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4,
      fft_q => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4,
      rd => logical2_y_net_x0,
      reset => logical1_y_net_x2,
      tx_reset => logical_y_net_x42,
      write => logical4_y_net_x1,
      i => reinterpret2_output_port_net_x1,
      occ => fifo_dcount_net_x3,
      q => reinterpret3_output_port_net_x1
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      clr => '0',
      ip(0) => delay2_q_net_x0,
      op(0) => inverter1_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      clr => '0',
      ip(0) => register2_q_net_x4,
      op(0) => inverter3_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x3,
      d1(0) => inverter1_op_net,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x3,
      d1(0) => convert2_dout_net_x4,
      d2(0) => register_q_net_x1,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net,
      d1(0) => register2_q_net_x4,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2,
      d1(0) => inverter3_op_net,
      y(0) => logical4_y_net_x1
    );

  mux: entity work.mux_bfe1d4f686
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      clr => '0',
      d0 => register2_q_net_x2,
      d1 => reinterpret2_output_port_net_x1,
      sel(0) => register1_q_net_x1,
      y => mux_y_net_x0
    );

  mux1: entity work.mux_bfe1d4f686
    port map (
      ce => ce_1_sg_x67,
      clk => clk_1_sg_x67,
      clr => '0',
      d0 => register3_q_net_x1,
      d1 => reinterpret3_output_port_net_x1,
      sel(0) => register1_q_net_x1,
      y => mux1_y_net_x1
    );

  posedge_35705d73cb: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      d => logical_y_net_x4,
      q => logical1_y_net_x2
    );

  preamble_gen_c25e867a97: entity work.preamble_gen_entity_c25e867a97
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      rd_en => convert2_dout_net_x4,
      tx_reset => logical_y_net_x42,
      tx_running => register2_q_net_x3,
      done => register1_q_net_x1,
      early_done => register_q_net_x1,
      i => register2_q_net_x2,
      q => register3_q_net_x1
    );

  relational1: entity work.relational_6dad3a03fc
    port map (
      a => fifo_dcount_net_x3,
      b(0) => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

  s_r_latch1_91a6112875: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      r => logical_y_net_x42,
      s => logical_y_net_x3,
      q => register2_q_net_x4
    );

  s_r_latch_c320bee3e4: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      r => logical_y_net_x42,
      s => logical1_y_net_x2,
      q => register2_q_net_x3
    );

  scaling_a269710a35: entity work.scaling_entity_a269710a35
    port map (
      ce_1 => ce_1_sg_x67,
      clk_1 => clk_1_sg_x67,
      i => mux_y_net_x0,
      preamble => delay1_q_net_x0,
      q => mux1_y_net_x1,
      regtx_scaling_payload => reinterpret1_output_port_net_x1,
      regtx_scaling_preamble => reinterpret_output_port_net_x1,
      i_x0 => mult_p_net_x1,
      q_x0 => mult1_p_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Registers/Status Bits"

entity status_bits_entity_a326423b7c is
  port (
    regtx_tx_running: in std_logic; 
    x32b: out std_logic_vector(31 downto 0)
  );
end status_bits_entity_a326423b7c;

architecture structural of status_bits_entity_a326423b7c is
  signal concat_y_net_x0: std_logic_vector(31 downto 0);
  signal constant_op_net: std_logic_vector(30 downto 0);
  signal register2_q_net_x0: std_logic;

begin
  register2_q_net_x0 <= regtx_tx_running;
  x32b <= concat_y_net_x0;

  concat: entity work.concat_e25f797841
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0 => constant_op_net,
      in1(0) => register2_q_net_x0,
      y => concat_y_net_x0
    );

  constant_x0: entity work.constant_bc7a810978
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Registers"

entity registers_entity_2d8965b1e5 is
  port (
    from_register1: in std_logic_vector(31 downto 0); 
    from_register2: in std_logic_vector(31 downto 0); 
    from_register3: in std_logic_vector(31 downto 0); 
    from_register4: in std_logic_vector(31 downto 0); 
    from_register5: in std_logic_vector(31 downto 0); 
    from_register6: in std_logic_vector(31 downto 0); 
    register2: in std_logic; 
    constant_x1: out std_logic; 
    regtx_anta_tx_en: out std_logic; 
    regtx_antb_tx_en: out std_logic; 
    regtx_cp_len: out std_logic_vector(7 downto 0); 
    regtx_fft_scaling: out std_logic_vector(5 downto 0); 
    regtx_num_sc: out std_logic_vector(7 downto 0); 
    regtx_pkt_buf_addr_offset: out std_logic_vector(7 downto 0); 
    regtx_pkt_buf_sel: out std_logic_vector(3 downto 0); 
    regtx_posttx_extension: out std_logic_vector(7 downto 0); 
    regtx_posttx_rf_en_extension: out std_logic_vector(7 downto 0); 
    regtx_posttx_rxsig_valid: out std_logic_vector(7 downto 0); 
    regtx_rc_rxen_enable: out std_logic; 
    regtx_reset: out std_logic; 
    regtx_reset_scrambling_lfsr_perpkt: out std_logic; 
    regtx_scaling_payload: out std_logic_vector(15 downto 0); 
    regtx_scaling_preamble: out std_logic_vector(15 downto 0); 
    regtx_start_direct: out std_logic; 
    regtx_start_indirect: out std_logic; 
    status_bits: out std_logic_vector(31 downto 0)
  );
end registers_entity_2d8965b1e5;

architecture structural of registers_entity_2d8965b1e5 is
  signal b_0_1_y_net_x0: std_logic;
  signal b_15_0_y_net: std_logic_vector(15 downto 0);
  signal b_15_8_1_y_net_x0: std_logic_vector(7 downto 0);
  signal b_15_8_y_net_x3: std_logic_vector(7 downto 0);
  signal b_1_y_net_x0: std_logic;
  signal b_1_y_net_x1: std_logic;
  signal b_23_16_y_net: std_logic_vector(7 downto 0);
  signal b_23_16_y_net_x2: std_logic_vector(7 downto 0);
  signal b_29_24_y_net_x1: std_logic_vector(5 downto 0);
  signal b_2_y_net_x1: std_logic;
  signal b_31_16_y_net: std_logic_vector(15 downto 0);
  signal b_31_y_net: std_logic;
  signal b_3_0_y_net: std_logic_vector(3 downto 0);
  signal b_3_y_net_x1: std_logic;
  signal b_7_0_1_y_net_x0: std_logic_vector(7 downto 0);
  signal b_7_0_y_net_x4: std_logic_vector(7 downto 0);
  signal concat_y_net_x1: std_logic_vector(31 downto 0);
  signal constant_op_net_x0: std_logic;
  signal from_register1_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register2_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register3_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register4_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register5_data_out_net_x0: std_logic_vector(31 downto 0);
  signal from_register6_data_out_net_x0: std_logic_vector(31 downto 0);
  signal lsb_y_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net_x2: std_logic_vector(15 downto 0);

begin
  from_register1_data_out_net_x0 <= from_register1;
  from_register2_data_out_net_x0 <= from_register2;
  from_register3_data_out_net_x0 <= from_register3;
  from_register4_data_out_net_x0 <= from_register4;
  from_register5_data_out_net_x0 <= from_register5;
  from_register6_data_out_net_x0 <= from_register6;
  register2_q_net_x1 <= register2;
  constant_x1 <= constant_op_net_x0;
  regtx_anta_tx_en <= b_2_y_net_x1;
  regtx_antb_tx_en <= b_3_y_net_x1;
  regtx_cp_len <= b_15_8_y_net_x3;
  regtx_fft_scaling <= b_29_24_y_net_x1;
  regtx_num_sc <= b_7_0_y_net_x4;
  regtx_pkt_buf_addr_offset <= b_23_16_y_net_x2;
  regtx_pkt_buf_sel <= b_3_0_y_net;
  regtx_posttx_extension <= b_7_0_1_y_net_x0;
  regtx_posttx_rf_en_extension <= b_15_8_1_y_net_x0;
  regtx_posttx_rxsig_valid <= b_23_16_y_net;
  regtx_rc_rxen_enable <= b_0_1_y_net_x0;
  regtx_reset <= b_31_y_net;
  regtx_reset_scrambling_lfsr_perpkt <= b_1_y_net_x0;
  regtx_scaling_payload <= reinterpret1_output_port_net_x2;
  regtx_scaling_preamble <= reinterpret_output_port_net_x2;
  regtx_start_direct <= lsb_y_net_x0;
  regtx_start_indirect <= b_1_y_net_x1;
  status_bits <= concat_y_net_x1;

  b_0_1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_0_1_y_net_x0
    );

  b_1: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_1_y_net_x0
    );

  b_15_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 15,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => from_register3_data_out_net_x0,
      y => b_15_0_y_net
    );

  b_15_8: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_15_8_y_net_x3
    );

  b_15_8_1: entity work.xlslice
    generic map (
      new_lsb => 8,
      new_msb => 15,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_15_8_1_y_net_x0
    );

  b_1_x0: entity work.xlslice
    generic map (
      new_lsb => 1,
      new_msb => 1,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register2_data_out_net_x0,
      y(0) => b_1_y_net_x1
    );

  b_2: entity work.xlslice
    generic map (
      new_lsb => 2,
      new_msb => 2,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_2_y_net_x1
    );

  b_23_16: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_23_16_y_net
    );

  b_23_16_x0: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 23,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register4_data_out_net_x0,
      y => b_23_16_y_net_x2
    );

  b_29_24: entity work.xlslice
    generic map (
      new_lsb => 24,
      new_msb => 29,
      x_width => 32,
      y_width => 6
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_29_24_y_net_x1
    );

  b_3: entity work.xlslice
    generic map (
      new_lsb => 3,
      new_msb => 3,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_3_y_net_x1
    );

  b_31: entity work.xlslice
    generic map (
      new_lsb => 31,
      new_msb => 31,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register5_data_out_net_x0,
      y(0) => b_31_y_net
    );

  b_31_16: entity work.xlslice
    generic map (
      new_lsb => 16,
      new_msb => 31,
      x_width => 32,
      y_width => 16
    )
    port map (
      x => from_register3_data_out_net_x0,
      y => b_31_16_y_net
    );

  b_3_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 3,
      x_width => 32,
      y_width => 4
    )
    port map (
      x => from_register4_data_out_net_x0,
      y => b_3_0_y_net
    );

  b_7_0: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register1_data_out_net_x0,
      y => b_7_0_y_net_x4
    );

  b_7_0_1: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 7,
      x_width => 32,
      y_width => 8
    )
    port map (
      x => from_register6_data_out_net_x0,
      y => b_7_0_1_y_net_x0
    );

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net_x0
    );

  lsb: entity work.xlslice
    generic map (
      new_lsb => 0,
      new_msb => 0,
      x_width => 32,
      y_width => 1
    )
    port map (
      x => from_register2_data_out_net_x0,
      y(0) => lsb_y_net_x0
    );

  reinterpret: entity work.reinterpret_ddc3ebdd7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => b_15_0_y_net,
      output_port => reinterpret_output_port_net_x2
    );

  reinterpret1: entity work.reinterpret_ddc3ebdd7c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      input_port => b_31_16_y_net,
      output_port => reinterpret1_output_port_net_x2
    );

  status_bits_a326423b7c: entity work.status_bits_entity_a326423b7c
    port map (
      regtx_tx_running => register2_q_net_x1,
      x32b => concat_y_net_x1
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Resets"

entity resets_entity_24d0a1b807 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    last_samp_output_to_dacs: in std_logic; 
    regtx_reset: in std_logic; 
    signal_decode_error: in std_logic; 
    tx_force_reset: out std_logic; 
    tx_phy_done: out std_logic; 
    tx_reset: out std_logic
  );
end resets_entity_24d0a1b807;

architecture structural of resets_entity_24d0a1b807 is
  signal b_31_y_net_x0: std_logic;
  signal ce_1_sg_x70: std_logic;
  signal clk_1_sg_x70: std_logic;
  signal constant_op_net: std_logic;
  signal convert1_dout_net_x0: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay_q_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical_y_net_x43: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register_q_net_x2: std_logic;
  signal simulation_multiplexer_dout_net: std_logic;

begin
  ce_1_sg_x70 <= ce_1;
  clk_1_sg_x70 <= clk_1;
  delay2_q_net_x1 <= last_samp_output_to_dacs;
  b_31_y_net_x0 <= regtx_reset;
  register_q_net_x2 <= signal_decode_error;
  tx_force_reset <= convert1_dout_net_x0;
  tx_phy_done <= logical1_y_net_x4;
  tx_reset <= logical_y_net_x43;

  constant_x0: entity work.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x70,
      clk => clk_1_sg_x70,
      clr => '0',
      din(0) => b_31_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net_x0
    );

  delay: entity work.xldelay
    generic map (
      latency => 16,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x70,
      clk => clk_1_sg_x70,
      d(0) => register2_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x0
    );

  logical: entity work.logical_6cb8f0ce02
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => simulation_multiplexer_dout_net,
      d1(0) => convert1_dout_net_x0,
      d2(0) => register2_q_net_x0,
      y(0) => logical_y_net_x43
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay2_q_net_x1,
      d1(0) => register_q_net_x2,
      y(0) => logical1_y_net_x1
    );

  posedge1_cd01046e00: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      d => logical1_y_net_x1,
      q => logical1_y_net_x4
    );

  s_r_latch_3226b7fe2e: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x70,
      clk_1 => clk_1_sg_x70,
      r => delay_q_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x0
    );

  simulation_multiplexer: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => constant_op_net,
      dout(0) => simulation_multiplexer_dout_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode/Conv Enc"

entity conv_enc_entity_0d273a2572 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    a: out std_logic; 
    b: out std_logic
  );
end conv_enc_entity_0d273a2572;

architecture structural of conv_enc_entity_0d273a2572 is
  signal a_xor_y_net_x0: std_logic;
  signal b_xor_y_net_x0: std_logic;
  signal ce_1_sg_x71: std_logic;
  signal clk_1_sg_x71: std_logic;
  signal convert2_dout_net: std_logic;
  signal convert_dout_net: std_logic;
  signal delay_q_net_x3: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x44: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x71 <= ce_1;
  clk_1_sg_x71 <= clk_1;
  logical_y_net_x0 <= data;
  delay_q_net_x3 <= en;
  logical_y_net_x44 <= rst;
  a <= a_xor_y_net_x0;
  b <= b_xor_y_net_x0;

  a_xor: entity work.logical_899cf9b568
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      d0(0) => logical_y_net_x0,
      d1(0) => register1_q_net,
      d2(0) => register2_q_net,
      d3(0) => register4_q_net,
      d4(0) => register5_q_net,
      en(0) => convert2_dout_net,
      y(0) => a_xor_y_net_x0
    );

  b_xor: entity work.logical_899cf9b568
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      d0(0) => logical_y_net_x0,
      d1(0) => register_q_net,
      d2(0) => register1_q_net,
      d3(0) => register2_q_net,
      d4(0) => register5_q_net,
      en(0) => convert2_dout_net,
      y(0) => b_xor_y_net_x0
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din(0) => logical_y_net_x44,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      clr => '0',
      din(0) => delay_q_net_x3,
      en => "1",
      dout(0) => convert2_dout_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => register_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => register1_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => register2_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => register3_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => register4_q_net,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x71,
      clk => clk_1_sg_x71,
      d(0) => logical_y_net_x0,
      en(0) => convert2_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode/Puncture/Rate 2/3"

entity x3_entity_c8f92e4f81 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    skip: out std_logic
  );
end x3_entity_c8f92e4f81;

architecture structural of x3_entity_c8f92e4f81 is
  signal ce_1_sg_x73: std_logic;
  signal clk_1_sg_x73: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal logical1_y_net_x0: std_logic;
  signal logical_y_net_x45: std_logic;
  signal relational_op_net_x0: std_logic;
  signal x0_3_op_net: std_logic_vector(1 downto 0);

begin
  ce_1_sg_x73 <= ce_1;
  clk_1_sg_x73 <= clk_1;
  logical1_y_net_x0 <= en;
  logical_y_net_x45 <= rst;
  skip <= relational_op_net_x0;

  constant1: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  relational: entity work.relational_5f1eb17108
    port map (
      a => x0_3_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net_x0
    );

  x0_3: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_6454489cfe866515",
      op_arith => xlUnsigned,
      op_width => 2
    )
    port map (
      ce => ce_1_sg_x73,
      clk => clk_1_sg_x73,
      clr => '0',
      en(0) => logical1_y_net_x0,
      rst(0) => logical_y_net_x45,
      op => x0_3_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode/Puncture/Rate 3/4"

entity x4_entity_1e2ac86547 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    rst: in std_logic; 
    skip: out std_logic
  );
end x4_entity_1e2ac86547;

architecture structural of x4_entity_1e2ac86547 is
  signal ce_1_sg_x74: std_logic;
  signal clk_1_sg_x74: std_logic;
  signal constant1_op_net: std_logic_vector(1 downto 0);
  signal constant2_op_net: std_logic_vector(2 downto 0);
  signal logical1_y_net_x1: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x46: std_logic;
  signal relational2_op_net: std_logic;
  signal relational_op_net: std_logic;
  signal x0_5_op_net: std_logic_vector(2 downto 0);

begin
  ce_1_sg_x74 <= ce_1;
  clk_1_sg_x74 <= clk_1;
  logical1_y_net_x1 <= en;
  logical_y_net_x46 <= rst;
  skip <= logical2_y_net_x0;

  constant1: entity work.constant_3a9a3daeb9
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant1_op_net
    );

  constant2: entity work.constant_469094441c
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational_op_net,
      d1(0) => relational2_op_net,
      y(0) => logical2_y_net_x0
    );

  relational: entity work.relational_706b9eb7ce
    port map (
      a => x0_5_op_net,
      b => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational2: entity work.relational_8fc7f5539b
    port map (
      a => x0_5_op_net,
      b => constant2_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational2_op_net
    );

  x0_5: entity work.xlcounter_limit_wlan_phy_tx_pmd
    generic map (
      cnt_15_0 => 5,
      cnt_31_16 => 0,
      cnt_47_32 => 0,
      cnt_63_48 => 0,
      core_name0 => "cntr_11_0_bcc28bfecf25caff",
      count_limited => 1,
      op_arith => xlUnsigned,
      op_width => 3
    )
    port map (
      ce => ce_1_sg_x74,
      clk => clk_1_sg_x74,
      clr => '0',
      en(0) => logical1_y_net_x1,
      rst(0) => logical_y_net_x46,
      op => x0_5_op_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode/Puncture"

entity puncture_entity_2dc0a9ab8c is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data: in std_logic; 
    data_bit_valid: in std_logic; 
    reset: in std_logic; 
    signal_code_rate: in std_logic_vector(1 downto 0); 
    coded_bit_tvalid: out std_logic
  );
end puncture_entity_2dc0a9ab8c;

architecture structural of puncture_entity_2dc0a9ab8c is
  signal ce_1_sg_x76: std_logic;
  signal clk_1_sg_x76: std_logic;
  signal concat_y_net: std_logic_vector(1 downto 0);
  signal convert1_dout_net: std_logic;
  signal convert6_dout_net_x2: std_logic_vector(1 downto 0);
  signal delay_q_net: std_logic;
  signal delay_q_net_x4: std_logic;
  signal inverter1_op_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical2_y_net: std_logic_vector(1 downto 0);
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net: std_logic;
  signal logical_y_net_x48: std_logic;
  signal mux1_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;
  signal relational_op_net_x0: std_logic;

begin
  ce_1_sg_x76 <= ce_1;
  clk_1_sg_x76 <= clk_1;
  logical1_y_net_x4 <= data;
  delay_q_net_x4 <= data_bit_valid;
  logical_y_net_x48 <= reset;
  convert6_dout_net_x2 <= signal_code_rate;
  coded_bit_tvalid <= mux1_y_net_x0;

  concat: entity work.concat_e6f5ee726b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      in0(0) => convert1_dout_net,
      in1(0) => convert1_dout_net,
      y => concat_y_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      din(0) => register2_q_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      d(0) => delay_q_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      ip(0) => relational_op_net_x0,
      op(0) => inverter_op_net
    );

  inverter1: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x76,
      clk => clk_1_sg_x76,
      clr => '0',
      ip(0) => logical2_y_net_x0,
      op(0) => inverter1_op_net
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x4,
      d1(0) => delay_q_net,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_33c9a0c803
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => concat_y_net,
      d1 => convert6_dout_net_x2,
      y => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => inverter_op_net,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => inverter1_op_net,
      y(0) => logical4_y_net
    );

  mux1: entity work.mux_472286caed
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x1,
      d1(0) => logical3_y_net,
      d2(0) => logical4_y_net,
      sel => logical2_y_net,
      y(0) => mux1_y_net_x0
    );

  posedge_fd5936ef1a: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      d => logical1_y_net_x4,
      q => logical1_y_net_x2
    );

  s_r_latch_d581cc219b: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      r => logical_y_net_x48,
      s => logical1_y_net_x2,
      q => register2_q_net_x0
    );

  x3_c8f92e4f81: entity work.x3_entity_c8f92e4f81
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      en => logical1_y_net_x1,
      rst => logical_y_net_x48,
      skip => relational_op_net_x0
    );

  x4_1e2ac86547: entity work.x4_entity_1e2ac86547
    port map (
      ce_1 => ce_1_sg_x76,
      clk_1 => clk_1_sg_x76,
      en => logical1_y_net_x1,
      rst => logical_y_net_x48,
      skip => logical2_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode/Scrambling LFSR"

entity scrambling_lfsr_entity_a68c54d78a is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    regtx_reset_scrambling_lfsr_perpkt: in std_logic; 
    tx_reset: in std_logic; 
    q: out std_logic
  );
end scrambling_lfsr_entity_a68c54d78a;

architecture structural of scrambling_lfsr_entity_a68c54d78a is
  signal assert1_dout_net: std_logic;
  signal assert_dout_net: std_logic;
  signal b_1_y_net_x1: std_logic;
  signal ce_1_sg_x77: std_logic;
  signal clk_1_sg_x77: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net: std_logic;
  signal logical_y_net_x49: std_logic;
  signal register1_q_net: std_logic;
  signal register2_q_net: std_logic;
  signal register3_q_net: std_logic;
  signal register4_q_net: std_logic;
  signal register5_q_net: std_logic;
  signal register6_q_net: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x77 <= ce_1;
  clk_1_sg_x77 <= clk_1;
  logical2_y_net_x0 <= en;
  b_1_y_net_x1 <= regtx_reset_scrambling_lfsr_perpkt;
  logical_y_net_x49 <= tx_reset;
  q <= convert2_dout_net_x0;

  assert1: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register3_q_net,
      dout(0) => assert1_dout_net
    );

  assert_x0: entity work.xlpassthrough
    generic map (
      din_width => 1,
      dout_width => 1
    )
    port map (
      din(0) => register6_q_net,
      dout(0) => assert_dout_net
    );

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      din(0) => logical1_y_net,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      din(0) => logical2_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      clr => '0',
      din(0) => logical_y_net,
      en => "1",
      dout(0) => convert2_dout_net_x0
    );

  logical: entity work.logical_e77c53f8bd
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => assert_dout_net,
      d1(0) => assert1_dout_net,
      y(0) => logical_y_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical_y_net_x49,
      d1(0) => b_1_y_net_x1,
      y(0) => logical1_y_net
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register1_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register2_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register3_q_net
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register3_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register4_q_net
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register4_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register5_q_net
    );

  register6: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => register5_q_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register6_q_net
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"1"
    )
    port map (
      ce => ce_1_sg_x77,
      clk => clk_1_sg_x77,
      d(0) => logical_y_net,
      en(0) => convert1_dout_net,
      rst(0) => convert_dout_net,
      q(0) => register_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Scramble & Encode"

entity \scramble___encode_entity_5f70e14e46\ is
  port (
    bit: in std_logic; 
    bit_source: in std_logic_vector(1 downto 0); 
    bit_valid: in std_logic; 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    data_pad_fcs: in std_logic; 
    registers: in std_logic; 
    tail: in std_logic; 
    tx_reset: in std_logic; 
    enc_bit: out std_logic; 
    enc_bit_valid: out std_logic
  );
end \scramble___encode_entity_5f70e14e46\;

architecture structural of \scramble___encode_entity_5f70e14e46\ is
  signal a_xor_y_net_x0: std_logic;
  signal b_1_y_net_x2: std_logic;
  signal b_xor_y_net_x0: std_logic;
  signal ce_1_sg_x78: std_logic;
  signal clk_1_sg_x78: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal convert2_dout_net_x0: std_logic;
  signal convert6_dout_net_x3: std_logic_vector(1 downto 0);
  signal delay1_q_net: std_logic;
  signal delay4_q_net_x1: std_logic;
  signal delay_q_net_x10: std_logic;
  signal delay_q_net_x5: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical_y_net_x0: std_logic;
  signal logical_y_net_x50: std_logic;
  signal mux1_y_net_x0: std_logic;
  signal mux_y_net_x7: std_logic;
  signal mux_y_net_x8: std_logic;

begin
  mux_y_net_x7 <= bit;
  convert6_dout_net_x3 <= bit_source;
  delay_q_net_x5 <= bit_valid;
  ce_1_sg_x78 <= ce_1;
  clk_1_sg_x78 <= clk_1;
  logical1_y_net_x5 <= data_pad_fcs;
  b_1_y_net_x2 <= registers;
  delay4_q_net_x1 <= tail;
  logical_y_net_x50 <= tx_reset;
  enc_bit <= mux_y_net_x8;
  enc_bit_valid <= delay_q_net_x10;

  conv_enc_0d273a2572: entity work.conv_enc_entity_0d273a2572
    port map (
      ce_1 => ce_1_sg_x78,
      clk_1 => clk_1_sg_x78,
      data => logical_y_net_x0,
      en => delay_q_net_x5,
      rst => logical_y_net_x50,
      a => a_xor_y_net_x0,
      b => b_xor_y_net_x0
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      din(0) => logical1_y_net_x5,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      din(0) => inverter_op_net,
      en => "1",
      dout(0) => convert2_dout_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      d(0) => mux1_y_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net_x10
    );

  delay1: entity work.xldelay
    generic map (
      latency => 2,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      d(0) => delay_q_net_x5,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x78,
      clk => clk_1_sg_x78,
      clr => '0',
      ip(0) => delay4_q_net_x1,
      op(0) => inverter_op_net
    );

  logical: entity work.logical_9d76333483
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => mux_y_net_x7,
      d1(0) => logical1_y_net,
      y(0) => logical_y_net_x0
    );

  logical1: entity work.logical_7b6bf7e572
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert1_dout_net,
      d1(0) => convert2_dout_net_x0,
      d2(0) => convert2_dout_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net_x5,
      d1(0) => logical1_y_net_x5,
      y(0) => logical2_y_net_x0
    );

  mux: entity work.mux_112ed141f4
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => a_xor_y_net_x0,
      d1(0) => b_xor_y_net_x0,
      sel(0) => delay1_q_net,
      y(0) => mux_y_net_x8
    );

  puncture_2dc0a9ab8c: entity work.puncture_entity_2dc0a9ab8c
    port map (
      ce_1 => ce_1_sg_x78,
      clk_1 => clk_1_sg_x78,
      data => logical1_y_net_x5,
      data_bit_valid => delay_q_net_x5,
      reset => logical_y_net_x50,
      signal_code_rate => convert6_dout_net_x3,
      coded_bit_tvalid => mux1_y_net_x0
    );

  scrambling_lfsr_a68c54d78a: entity work.scrambling_lfsr_entity_a68c54d78a
    port map (
      ce_1 => ce_1_sg_x78,
      clk_1 => clk_1_sg_x78,
      en => logical2_y_net_x0,
      regtx_reset_scrambling_lfsr_perpkt => b_1_y_net_x2,
      tx_reset => logical_y_net_x50,
      q => convert2_dout_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Add Extension"

entity add_extension_entity_08b6a45d51 is
  port (
    ce_1: in std_logic; 
    ce_8: in std_logic; 
    clk_1: in std_logic; 
    clk_8: in std_logic; 
    iq_done: in std_logic; 
    regtx_posttx_extension: in std_logic_vector(7 downto 0); 
    rst: in std_logic; 
    tx_start: in std_logic; 
    tx_active: out std_logic
  );
end add_extension_entity_08b6a45d51;

architecture structural of add_extension_entity_08b6a45d51 is
  signal b_7_0_1_y_net_x1: std_logic_vector(7 downto 0);
  signal ce_1_sg_x81: std_logic;
  signal ce_8_sg_x0: std_logic;
  signal clk_1_sg_x81: std_logic;
  signal clk_8_sg_x0: std_logic;
  signal constant_op_net: std_logic;
  signal convert1_dout_net_x1: std_logic;
  signal counter1_op_net: std_logic_vector(7 downto 0);
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical2_y_net_x1: std_logic;
  signal logical_y_net_x6: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x2: std_logic;
  signal relational3_op_net: std_logic;
  signal up_sample_q_net: std_logic;

begin
  ce_1_sg_x81 <= ce_1;
  ce_8_sg_x0 <= ce_8;
  clk_1_sg_x81 <= clk_1;
  clk_8_sg_x0 <= clk_8;
  logical1_y_net_x6 <= iq_done;
  b_7_0_1_y_net_x1 <= regtx_posttx_extension;
  convert1_dout_net_x1 <= rst;
  logical_y_net_x6 <= tx_start;
  tx_active <= register2_q_net_x2;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_86806e294f737f4c",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x81,
      clk => clk_1_sg_x81,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => logical2_y_net_x1,
      op => counter1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => up_sample_q_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational3_op_net,
      d1(0) => convert1_dout_net_x1,
      y(0) => logical2_y_net_x1
    );

  relational3: entity work.relational_7bfd319389
    port map (
      a => counter1_op_net,
      b => b_7_0_1_y_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_65222083f7: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x81,
      clk_1 => clk_1_sg_x81,
      r => logical2_y_net_x1,
      s => logical1_y_net_x6,
      q => register2_q_net_x0
    );

  s_r_latch2_1b9d9de144: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x81,
      clk_1 => clk_1_sg_x81,
      r => logical2_y_net_x1,
      s => logical_y_net_x6,
      q => register2_q_net_x2
    );

  up_sample: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => constant_op_net,
      dest_ce => ce_1_sg_x81,
      dest_clk => clk_1_sg_x81,
      dest_clr => '0',
      en => "1",
      src_ce => ce_8_sg_x0,
      src_clk => clk_8_sg_x0,
      src_clr => '0',
      q(0) => up_sample_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Add Extension1"

entity add_extension1_entity_77211131cc is
  port (
    ce_1: in std_logic; 
    ce_8: in std_logic; 
    clk_1: in std_logic; 
    clk_8: in std_logic; 
    last_samp: in std_logic; 
    regtx_posttx_rf_en_extension: in std_logic_vector(7 downto 0); 
    regtx_posttx_rxsig_valid: in std_logic_vector(7 downto 0); 
    rst: in std_logic; 
    disable_rf_tx: out std_logic; 
    rxsig_valid: out std_logic
  );
end add_extension1_entity_77211131cc;

architecture structural of add_extension1_entity_77211131cc is
  signal b_15_8_1_y_net_x1: std_logic_vector(7 downto 0);
  signal b_23_16_y_net_x0: std_logic_vector(7 downto 0);
  signal ce_1_sg_x86: std_logic;
  signal ce_8_sg_x1: std_logic;
  signal clk_1_sg_x86: std_logic;
  signal clk_8_sg_x1: std_logic;
  signal constant_op_net: std_logic;
  signal convert1_dout_net_x2: std_logic;
  signal counter1_op_net: std_logic_vector(7 downto 0);
  signal logical1_y_net: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x10: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x9: std_logic;
  signal logical2_y_net_x0: std_logic;
  signal logical3_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;
  signal relational1_op_net_x0: std_logic;
  signal relational3_op_net: std_logic;
  signal up_sample_q_net: std_logic;

begin
  ce_1_sg_x86 <= ce_1;
  ce_8_sg_x1 <= ce_8;
  clk_1_sg_x86 <= clk_1;
  clk_8_sg_x1 <= clk_8;
  logical1_y_net_x9 <= last_samp;
  b_15_8_1_y_net_x1 <= regtx_posttx_rf_en_extension;
  b_23_16_y_net_x0 <= regtx_posttx_rxsig_valid;
  convert1_dout_net_x2 <= rst;
  disable_rf_tx <= logical1_y_net_x10;
  rxsig_valid <= logical1_y_net_x11;

  constant_x0: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant_op_net
    );

  counter1: entity work.xlcounter_free_wlan_phy_tx_pmd
    generic map (
      core_name0 => "cntr_11_0_86806e294f737f4c",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x86,
      clk => clk_1_sg_x86,
      clr => '0',
      en(0) => logical1_y_net,
      rst(0) => logical2_y_net_x0,
      op => counter1_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => register2_q_net_x0,
      d1(0) => up_sample_q_net,
      y(0) => logical1_y_net
    );

  logical2: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x0,
      d1(0) => convert1_dout_net_x2,
      y(0) => logical2_y_net_x0
    );

  logical3: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational1_op_net_x0,
      d1(0) => relational3_op_net,
      y(0) => logical3_y_net_x0
    );

  posedge1_92e29d3358: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x86,
      clk_1 => clk_1_sg_x86,
      d => logical1_y_net_x9,
      q => logical1_y_net_x1
    );

  posedge2_38d01180e9: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x86,
      clk_1 => clk_1_sg_x86,
      d => logical3_y_net_x0,
      q => logical1_y_net_x10
    );

  posedge3_213ec870de: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x86,
      clk_1 => clk_1_sg_x86,
      d => relational1_op_net_x0,
      q => logical1_y_net_x11
    );

  relational1: entity work.relational_7bfd319389
    port map (
      a => counter1_op_net,
      b => b_23_16_y_net_x0,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net_x0
    );

  relational3: entity work.relational_7bfd319389
    port map (
      a => counter1_op_net,
      b => b_15_8_1_y_net_x1,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational3_op_net
    );

  s_r_latch1_45f12eaae9: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x86,
      clk_1 => clk_1_sg_x86,
      r => logical2_y_net_x0,
      s => logical1_y_net_x1,
      q => register2_q_net_x0
    );

  up_sample: entity work.xlusamp
    generic map (
      copy_samples => 0,
      d_arith => xlUnsigned,
      d_bin_pt => 0,
      d_width => 1,
      latency => 0,
      q_arith => xlUnsigned,
      q_bin_pt => 0,
      q_width => 1
    )
    port map (
      d(0) => constant_op_net,
      dest_ce => ce_1_sg_x86,
      dest_clk => clk_1_sg_x86,
      dest_clr => '0',
      en => "1",
      src_ce => ce_8_sg_x1,
      src_clk => clk_8_sg_x1,
      src_clr => '0',
      q(0) => up_sample_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/Pkt Buf Sel"

entity pkt_buf_sel_entity_412d479839 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    hw_tx: in std_logic; 
    phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    regtx_pkt_buf_sel: in std_logic_vector(3 downto 0); 
    sw_tx: in std_logic; 
    pkt_buf: out std_logic_vector(3 downto 0)
  );
end pkt_buf_sel_entity_412d479839;

architecture structural of pkt_buf_sel_entity_412d479839 is
  signal b_3_0_y_net_x0: std_logic_vector(3 downto 0);
  signal ce_1_sg_x87: std_logic;
  signal clk_1_sg_x87: std_logic;
  signal convert1_dout_net_x0: std_logic;
  signal convert1_dout_net_x1: std_logic;
  signal convert_dout_net: std_logic;
  signal logical1_y_net: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal mux_y_net_x2: std_logic_vector(3 downto 0);
  signal phy_tx_pkt_buf_net_x0: std_logic_vector(3 downto 0);
  signal register1_q_net: std_logic_vector(3 downto 0);
  signal register2_q_net: std_logic_vector(3 downto 0);
  signal register3_q_net: std_logic;

begin
  ce_1_sg_x87 <= ce_1;
  clk_1_sg_x87 <= clk_1;
  convert1_dout_net_x1 <= hw_tx;
  phy_tx_pkt_buf_net_x0 <= phy_tx_pkt_buf;
  b_3_0_y_net_x0 <= regtx_pkt_buf_sel;
  logical5_y_net_x0 <= sw_tx;
  pkt_buf <= mux_y_net_x2;

  convert: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      din(0) => logical5_y_net_x0,
      en => "1",
      dout(0) => convert_dout_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      clr => '0',
      din(0) => convert1_dout_net_x1,
      en => "1",
      dout(0) => convert1_dout_net_x0
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert_dout_net,
      d1(0) => convert1_dout_net_x0,
      y(0) => logical1_y_net
    );

  mux: entity work.mux_f9c0f11a18
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register1_q_net,
      d1 => register2_q_net,
      sel(0) => register3_q_net,
      y => mux_y_net_x2
    );

  register1: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      d => b_3_0_y_net_x0,
      en(0) => convert_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 4,
      init_value => b"0000"
    )
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      d => phy_tx_pkt_buf_net_x0,
      en(0) => convert1_dout_net_x0,
      rst => "0",
      q => register2_q_net
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x87,
      clk => clk_1_sg_x87,
      d(0) => convert1_dout_net_x0,
      en(0) => logical1_y_net,
      rst => "0",
      q(0) => register3_q_net
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/S-R Latch2"

entity s_r_latch2_entity_c31d9fc389 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    r: in std_logic; 
    s: in std_logic; 
    q: out std_logic
  );
end s_r_latch2_entity_c31d9fc389;

architecture structural of s_r_latch2_entity_c31d9fc389 is
  signal ce_1_sg_x94: std_logic;
  signal clk_1_sg_x94: std_logic;
  signal constant1_op_net: std_logic;
  signal convert1_dout_net: std_logic;
  signal convert2_dout_net: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;

begin
  ce_1_sg_x94 <= ce_1;
  clk_1_sg_x94 <= clk_1;
  logical8_y_net_x0 <= r;
  logical1_y_net_x4 <= s;
  q <= register2_q_net_x0;

  constant1: entity work.constant_6293007044
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      clr => '0',
      din(0) => logical8_y_net_x0,
      en => "1",
      dout(0) => convert1_dout_net
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      clr => '0',
      din(0) => logical1_y_net_x4,
      en => "1",
      dout(0) => convert2_dout_net
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x94,
      clk => clk_1_sg_x94,
      d(0) => constant1_op_net,
      en(0) => convert2_dout_net,
      rst(0) => convert1_dout_net,
      q(0) => register2_q_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/negedge"

entity negedge_entity_5ee9de3524 is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end negedge_entity_5ee9de3524;

architecture structural of negedge_entity_5ee9de3524 is
  signal ce_1_sg_x95: std_logic;
  signal clk_1_sg_x95: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal register2_q_net_x4: std_logic;

begin
  ce_1_sg_x95 <= ce_1;
  clk_1_sg_x95 <= clk_1;
  register2_q_net_x4 <= d;
  q <= logical1_y_net_x0;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      d(0) => register2_q_net_x4,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x95,
      clk => clk_1_sg_x95,
      clr => '0',
      ip(0) => register2_q_net_x4,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl/negedge1"

entity negedge1_entity_64a346f30b is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    d: in std_logic; 
    q: out std_logic
  );
end negedge1_entity_64a346f30b;

architecture structural of negedge1_entity_64a346f30b is
  signal ce_1_sg_x96: std_logic;
  signal clk_1_sg_x96: std_logic;
  signal delay_q_net: std_logic;
  signal inverter_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal register3_q_net_x0: std_logic;

begin
  ce_1_sg_x96 <= ce_1;
  clk_1_sg_x96 <= clk_1;
  register3_q_net_x0 <= d;
  q <= logical1_y_net_x0;

  delay: entity work.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      d(0) => register3_q_net_x0,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  inverter: entity work.inverter_e2b989a05e
    port map (
      ce => ce_1_sg_x96,
      clk => clk_1_sg_x96,
      clr => '0',
      ip(0) => register3_q_net_x0,
      op(0) => inverter_op_net
    );

  logical1: entity work.logical_938d99ac11
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => delay_q_net,
      d1(0) => inverter_op_net,
      y(0) => logical1_y_net_x0
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd/Start Ctrl"

entity start_ctrl_entity_3ba2a032ad is
  port (
    ce_1: in std_logic; 
    ce_8: in std_logic; 
    clk_1: in std_logic; 
    clk_8: in std_logic; 
    dac_tx_clk: in std_logic; 
    phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    phy_tx_start: in std_logic; 
    rc_phy_start: in std_logic; 
    registers: in std_logic_vector(7 downto 0); 
    registers_x0: in std_logic_vector(7 downto 0); 
    registers_x1: in std_logic_vector(3 downto 0); 
    registers_x2: in std_logic_vector(7 downto 0); 
    regtx_rc_rxen_enable: in std_logic; 
    regtx_start_direct: in std_logic; 
    regtx_start_indirect: in std_logic; 
    tx_force_reset: in std_logic; 
    tx_phy_done: in std_logic; 
    negedge_x0: out std_logic; 
    phy_start: out std_logic; 
    posedge2: out std_logic; 
    register1_x0: out std_logic; 
    register2_x0: out std_logic; 
    register4_x0: out std_logic; 
    register5_x0: out std_logic; 
    regtx_tx_running: out std_logic; 
    tx_iq_samp_ce: out std_logic; 
    tx_pkt_buf_sel: out std_logic_vector(3 downto 0)
  );
end start_ctrl_entity_3ba2a032ad;

architecture structural of start_ctrl_entity_3ba2a032ad is
  signal b_0_1_y_net_x1: std_logic;
  signal b_15_8_1_y_net_x2: std_logic_vector(7 downto 0);
  signal b_1_y_net_x2: std_logic;
  signal b_23_16_y_net_x1: std_logic_vector(7 downto 0);
  signal b_3_0_y_net_x1: std_logic_vector(3 downto 0);
  signal b_7_0_1_y_net_x2: std_logic_vector(7 downto 0);
  signal ce_1_sg_x97: std_logic;
  signal ce_8_sg_x2: std_logic;
  signal clk_1_sg_x97: std_logic;
  signal clk_8_sg_x2: std_logic;
  signal convert1_dout_net_x1: std_logic;
  signal convert1_dout_net_x3: std_logic;
  signal convert2_dout_net_x5: std_logic;
  signal convert3_dout_net: std_logic;
  signal convert4_dout_net_x0: std_logic;
  signal convert5_dout_net: std_logic;
  signal convert6_dout_net: std_logic;
  signal convert7_dout_net: std_logic;
  signal convert8_dout_net: std_logic;
  signal dac_tx_clk_net_x0: std_logic;
  signal delay1_q_net: std_logic;
  signal delay_q_net: std_logic;
  signal inverter2_op_net: std_logic;
  signal inverter3_op_net: std_logic;
  signal logical1_y_net_x0: std_logic;
  signal logical1_y_net_x1: std_logic;
  signal logical1_y_net_x11: std_logic;
  signal logical1_y_net_x12: std_logic;
  signal logical1_y_net_x13: std_logic;
  signal logical1_y_net_x14: std_logic;
  signal logical1_y_net_x15: std_logic;
  signal logical1_y_net_x3: std_logic;
  signal logical1_y_net_x4: std_logic;
  signal logical1_y_net_x6: std_logic;
  signal logical2_y_net: std_logic;
  signal logical3_y_net: std_logic;
  signal logical4_y_net_x0: std_logic;
  signal logical5_y_net_x0: std_logic;
  signal logical6_y_net_x0: std_logic;
  signal logical7_y_net_x0: std_logic;
  signal logical8_y_net_x0: std_logic;
  signal logical_y_net_x7: std_logic;
  signal lsb_y_net_x1: std_logic;
  signal mux_y_net_x3: std_logic_vector(3 downto 0);
  signal phy_tx_pkt_buf_net_x1: std_logic_vector(3 downto 0);
  signal phy_tx_start_net_x0: std_logic;
  signal rc_phy_start_net_x0: std_logic;
  signal register1_q_net_x0: std_logic;
  signal register2_q_net_x0: std_logic;
  signal register2_q_net_x1: std_logic;
  signal register2_q_net_x3: std_logic;
  signal register2_q_net_x4: std_logic;
  signal register2_q_net_x5: std_logic;
  signal register3_q_net_x0: std_logic;
  signal register4_q_net_x0: std_logic;
  signal register5_q_net_x0: std_logic;
  signal register_q_net: std_logic;

begin
  ce_1_sg_x97 <= ce_1;
  ce_8_sg_x2 <= ce_8;
  clk_1_sg_x97 <= clk_1;
  clk_8_sg_x2 <= clk_8;
  dac_tx_clk_net_x0 <= dac_tx_clk;
  phy_tx_pkt_buf_net_x1 <= phy_tx_pkt_buf;
  phy_tx_start_net_x0 <= phy_tx_start;
  rc_phy_start_net_x0 <= rc_phy_start;
  b_15_8_1_y_net_x2 <= registers;
  b_23_16_y_net_x1 <= registers_x0;
  b_3_0_y_net_x1 <= registers_x1;
  b_7_0_1_y_net_x2 <= registers_x2;
  b_0_1_y_net_x1 <= regtx_rc_rxen_enable;
  lsb_y_net_x1 <= regtx_start_direct;
  b_1_y_net_x2 <= regtx_start_indirect;
  convert1_dout_net_x3 <= tx_force_reset;
  logical1_y_net_x13 <= tx_phy_done;
  negedge_x0 <= logical1_y_net_x15;
  phy_start <= logical_y_net_x7;
  posedge2 <= logical1_y_net_x14;
  register1_x0 <= register1_q_net_x0;
  register2_x0 <= register2_q_net_x3;
  register4_x0 <= register4_q_net_x0;
  register5_x0 <= register5_q_net_x0;
  regtx_tx_running <= register2_q_net_x5;
  tx_iq_samp_ce <= convert2_dout_net_x5;
  tx_pkt_buf_sel <= mux_y_net_x3;

  add_extension1_77211131cc: entity work.add_extension1_entity_77211131cc
    port map (
      ce_1 => ce_1_sg_x97,
      ce_8 => ce_8_sg_x2,
      clk_1 => clk_1_sg_x97,
      clk_8 => clk_8_sg_x2,
      last_samp => logical1_y_net_x13,
      regtx_posttx_rf_en_extension => b_15_8_1_y_net_x2,
      regtx_posttx_rxsig_valid => b_23_16_y_net_x1,
      rst => convert1_dout_net_x3,
      disable_rf_tx => logical1_y_net_x11,
      rxsig_valid => logical1_y_net_x12
    );

  add_extension_08b6a45d51: entity work.add_extension_entity_08b6a45d51
    port map (
      ce_1 => ce_1_sg_x97,
      ce_8 => ce_8_sg_x2,
      clk_1 => clk_1_sg_x97,
      clk_8 => clk_8_sg_x2,
      iq_done => logical1_y_net_x13,
      regtx_posttx_extension => b_7_0_1_y_net_x2,
      rst => convert1_dout_net_x3,
      tx_start => logical_y_net_x7,
      tx_active => register2_q_net_x4
    );

  convert1: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => phy_tx_start_net_x0,
      en => "1",
      dout(0) => convert1_dout_net_x1
    );

  convert2: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => logical1_y_net_x6,
      en => "1",
      dout(0) => convert2_dout_net_x5
    );

  convert3: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => b_1_y_net_x2,
      en => "1",
      dout(0) => convert3_dout_net
    );

  convert4: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => b_0_1_y_net_x1,
      en => "1",
      dout(0) => convert4_dout_net_x0
    );

  convert5: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => lsb_y_net_x1,
      en => "1",
      dout(0) => convert5_dout_net
    );

  convert6: entity work.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => rc_phy_start_net_x0,
      en => "1",
      dout(0) => convert6_dout_net
    );

  convert7: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => logical2_y_net,
      en => "1",
      dout(0) => convert7_dout_net
    );

  convert8: entity work.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      din(0) => logical3_y_net,
      en => "1",
      dout(0) => convert8_dout_net
    );

  delay: entity work.xldelay
    generic map (
      latency => 32,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => logical2_y_net,
      en => '1',
      rst => '1',
      q(0) => delay_q_net
    );

  delay1: entity work.xldelay
    generic map (
      latency => 32,
      reg_retiming => 0,
      reset => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => logical3_y_net,
      en => '1',
      rst => '1',
      q(0) => delay1_q_net
    );

  inverter2: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      ip(0) => delay_q_net,
      op(0) => inverter2_op_net
    );

  inverter3: entity work.inverter_e5b38cca3b
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      clr => '0',
      ip(0) => delay1_q_net,
      op(0) => inverter3_op_net
    );

  logical: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert5_dout_net,
      d1(0) => convert6_dout_net,
      y(0) => logical_y_net_x7
    );

  logical1: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert3_dout_net,
      d1(0) => convert1_dout_net_x1,
      y(0) => logical1_y_net_x1
    );

  logical2: entity work.logical_954ee29728
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert4_dout_net_x0,
      d1(0) => register2_q_net_x0,
      d2(0) => inverter3_op_net,
      y(0) => logical2_y_net
    );

  logical3: entity work.logical_80f90b97d0
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => inverter2_op_net,
      d1(0) => register2_q_net_x5,
      y(0) => logical3_y_net
    );

  logical4: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x0,
      d1(0) => logical1_y_net_x3,
      y(0) => logical4_y_net_x0
    );

  logical5: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => convert3_dout_net,
      d1(0) => convert5_dout_net,
      y(0) => logical5_y_net_x0
    );

  logical6: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical4_y_net_x0,
      d1(0) => convert1_dout_net_x3,
      y(0) => logical6_y_net_x0
    );

  logical7: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x4,
      d1(0) => convert1_dout_net_x3,
      y(0) => logical7_y_net_x0
    );

  logical8: entity work.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => logical1_y_net_x12,
      d1(0) => convert1_dout_net_x3,
      y(0) => logical8_y_net_x0
    );

  negedge1_64a346f30b: entity work.negedge1_entity_64a346f30b
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => register3_q_net_x0,
      q => logical1_y_net_x6
    );

  negedge_5ee9de3524: entity work.negedge_entity_5ee9de3524
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => register2_q_net_x4,
      q => logical1_y_net_x15
    );

  pkt_buf_sel_412d479839: entity work.pkt_buf_sel_entity_412d479839
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      hw_tx => convert1_dout_net_x1,
      phy_tx_pkt_buf => phy_tx_pkt_buf_net_x1,
      regtx_pkt_buf_sel => b_3_0_y_net_x1,
      sw_tx => logical5_y_net_x0,
      pkt_buf => mux_y_net_x3
    );

  posedge1_95d3e0d45f: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => logical1_y_net_x1,
      q => logical1_y_net_x4
    );

  posedge2_6c78090f16: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => register2_q_net_x4,
      q => logical1_y_net_x14
    );

  posedge3_52a7b75f24: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => logical1_y_net_x11,
      q => logical1_y_net_x3
    );

  posedge_ebc0a6d5d0: entity work.posedge1_entity_9966c21e4f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      d => convert4_dout_net_x0,
      q => logical1_y_net_x0
    );

  register1: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => register_q_net,
      en => "1",
      rst => "0",
      q(0) => register1_q_net_x0
    );

  register2: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => register2_q_net_x1,
      en => "1",
      rst => "0",
      q(0) => register2_q_net_x3
    );

  register3: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => dac_tx_clk_net_x0,
      en => "1",
      rst => "0",
      q(0) => register3_q_net_x0
    );

  register4: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => convert7_dout_net,
      en => "1",
      rst => "0",
      q(0) => register4_q_net_x0
    );

  register5: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => convert8_dout_net,
      en => "1",
      rst => "0",
      q(0) => register5_q_net_x0
    );

  register_x0: entity work.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x97,
      clk => clk_1_sg_x97,
      d(0) => register2_q_net_x4,
      en => "1",
      rst => "0",
      q(0) => register_q_net
    );

  s_r_latch1_96bb620271: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      r => logical7_y_net_x0,
      s => logical4_y_net_x0,
      q => register2_q_net_x0
    );

  s_r_latch2_c31d9fc389: entity work.s_r_latch2_entity_c31d9fc389
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      r => logical8_y_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x1
    );

  s_r_latch_9c9835a519: entity work.s_r_latch1_entity_7106e36b8f
    port map (
      ce_1 => ce_1_sg_x97,
      clk_1 => clk_1_sg_x97,
      r => logical6_y_net_x0,
      s => logical1_y_net_x4,
      q => register2_q_net_x5
    );

end structural;
library IEEE;
use IEEE.std_logic_1164.all;
use work.conv_pkg.all;

-- Generated from Simulink block "wlan_phy_tx_pmd"

entity wlan_phy_tx_pmd is
  port (
    axi_aresetn: in std_logic; 
    bram_din: in std_logic_vector(63 downto 0); 
    ce_1: in std_logic; 
    ce_8: in std_logic; 
    clk_1: in std_logic; 
    clk_8: in std_logic; 
    dac_tx_clk: in std_logic; 
    data_out: in std_logic_vector(31 downto 0); 
    data_out_x0: in std_logic_vector(31 downto 0); 
    data_out_x1: in std_logic_vector(31 downto 0); 
    data_out_x2: in std_logic_vector(31 downto 0); 
    data_out_x3: in std_logic_vector(31 downto 0); 
    data_out_x4: in std_logic_vector(31 downto 0); 
    data_out_x5: in std_logic_vector(31 downto 0); 
    dout: in std_logic_vector(31 downto 0); 
    dout_x0: in std_logic_vector(31 downto 0); 
    dout_x1: in std_logic_vector(31 downto 0); 
    dout_x2: in std_logic_vector(31 downto 0); 
    dout_x3: in std_logic_vector(31 downto 0); 
    dout_x4: in std_logic_vector(31 downto 0); 
    phy_tx_pkt_buf: in std_logic_vector(3 downto 0); 
    phy_tx_start: in std_logic; 
    plb_ce_1: in std_logic; 
    plb_clk_1: in std_logic; 
    rc_phy_start: in std_logic; 
    s_axi_araddr: in std_logic_vector(31 downto 0); 
    s_axi_arburst: in std_logic_vector(1 downto 0); 
    s_axi_arcache: in std_logic_vector(3 downto 0); 
    s_axi_arid: in std_logic_vector(7 downto 0); 
    s_axi_arlen: in std_logic_vector(7 downto 0); 
    s_axi_arlock: in std_logic_vector(1 downto 0); 
    s_axi_arprot: in std_logic_vector(2 downto 0); 
    s_axi_arsize: in std_logic_vector(2 downto 0); 
    s_axi_arvalid: in std_logic; 
    s_axi_awaddr: in std_logic_vector(31 downto 0); 
    s_axi_awburst: in std_logic_vector(1 downto 0); 
    s_axi_awcache: in std_logic_vector(3 downto 0); 
    s_axi_awid: in std_logic_vector(7 downto 0); 
    s_axi_awlen: in std_logic_vector(7 downto 0); 
    s_axi_awlock: in std_logic_vector(1 downto 0); 
    s_axi_awprot: in std_logic_vector(2 downto 0); 
    s_axi_awsize: in std_logic_vector(2 downto 0); 
    s_axi_awvalid: in std_logic; 
    s_axi_bready: in std_logic; 
    s_axi_rready: in std_logic; 
    s_axi_wdata: in std_logic_vector(31 downto 0); 
    s_axi_wlast: in std_logic; 
    s_axi_wstrb: in std_logic_vector(3 downto 0); 
    s_axi_wvalid: in std_logic; 
    bram_addr: out std_logic_vector(31 downto 0); 
    bram_dout: out std_logic_vector(63 downto 0); 
    bram_en: out std_logic; 
    bram_reset: out std_logic; 
    bram_wen: out std_logic_vector(7 downto 0); 
    data_in: out std_logic_vector(31 downto 0); 
    data_in_x0: out std_logic_vector(31 downto 0); 
    data_in_x1: out std_logic_vector(31 downto 0); 
    data_in_x2: out std_logic_vector(31 downto 0); 
    data_in_x3: out std_logic_vector(31 downto 0); 
    data_in_x4: out std_logic_vector(31 downto 0); 
    data_in_x5: out std_logic_vector(31 downto 0); 
    dbg_tx_running: out std_logic; 
    en: out std_logic; 
    en_x0: out std_logic; 
    en_x1: out std_logic; 
    en_x2: out std_logic; 
    en_x3: out std_logic; 
    en_x4: out std_logic; 
    en_x5: out std_logic; 
    phy_tx_done: out std_logic; 
    phy_tx_started: out std_logic; 
    rc_usr_rxen: out std_logic; 
    rc_usr_txen: out std_logic; 
    rfa_dac_i: out std_logic_vector(11 downto 0); 
    rfa_dac_q: out std_logic_vector(11 downto 0); 
    rfb_dac_i: out std_logic_vector(11 downto 0); 
    rfb_dac_q: out std_logic_vector(11 downto 0); 
    rx_sigs_invalid: out std_logic; 
    s_axi_arready: out std_logic; 
    s_axi_awready: out std_logic; 
    s_axi_bid: out std_logic_vector(7 downto 0); 
    s_axi_bresp: out std_logic_vector(1 downto 0); 
    s_axi_bvalid: out std_logic; 
    s_axi_rdata: out std_logic_vector(31 downto 0); 
    s_axi_rid: out std_logic_vector(7 downto 0); 
    s_axi_rlast: out std_logic; 
    s_axi_rresp: out std_logic_vector(1 downto 0); 
    s_axi_rvalid: out std_logic; 
    s_axi_wready: out std_logic
  );
end wlan_phy_tx_pmd;

architecture structural of wlan_phy_tx_pmd is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "wlan_phy_tx_pmd,sysgen_core,{clock_period=6.25000000,clocking=Clock_Enables,sample_periods=1.00000000000 8.00000000000 1.00000000000,testbench=0,total_blocks=1810,xilinx_accumulator_block=1,xilinx_adder_subtracter_block=5,xilinx_arithmetic_relational_operator_block=35,xilinx_assert_block=12,xilinx_axi_fifo_block_block=1,xilinx_bit_slice_extractor_block=110,xilinx_bus_concatenator_block=26,xilinx_bus_multiplexer_block=27,xilinx_constant_block_block=111,xilinx_counter_block=15,xilinx_delay_block=68,xilinx_disregard_subsystem_for_generation_block=2,xilinx_dual_port_random_access_memory_block=4,xilinx_edk_core_block=1,xilinx_edk_processor_block=1,xilinx_fast_fourier_transform_8_0__block=1,xilinx_fifo_block_block=1,xilinx_gateway_in_block=31,xilinx_gateway_out_block=203,xilinx_inverter_block=57,xilinx_logical_block_block=112,xilinx_mcode_block_block=1,xilinx_multiplier_block=2,xilinx_register_block=67,xilinx_shared_memory_based_from_register_block=7,xilinx_shared_memory_based_to_register_block=7,xilinx_simulation_multiplexer_block=2,xilinx_single_port_read_only_memory_block=10,xilinx_system_generator_block=1,xilinx_type_converter_block=91,xilinx_type_reinterpreter_block=11,xilinx_up_sampler_block=2,}";

  signal axi_aresetn_net: std_logic;
  signal axi_fifo_m_axis_tvalid_net_x2: std_logic;
  signal axi_fifo_s_axis_tready_net_x2: std_logic;
  signal b_0_1_y_net_x1: std_logic;
  signal b_15_8_1_y_net_x2: std_logic_vector(7 downto 0);
  signal b_15_8_y_net_x3: std_logic_vector(7 downto 0);
  signal b_1_y_net_x2: std_logic;
  signal b_1_y_net_x3: std_logic;
  signal b_23_16_y_net_x1: std_logic_vector(7 downto 0);
  signal b_23_16_y_net_x2: std_logic_vector(7 downto 0);
  signal b_29_24_y_net_x1: std_logic_vector(5 downto 0);
  signal b_2_1_y_net_x1: std_logic_vector(1 downto 0);
  signal b_2_y_net_x1: std_logic;
  signal b_31_y_net_x0: std_logic;
  signal b_3_0_y_net_x1: std_logic_vector(3 downto 0);
  signal b_3_y_net_x1: std_logic;
  signal b_7_0_1_y_net_x2: std_logic_vector(7 downto 0);
  signal b_7_0_y_net_x4: std_logic_vector(7 downto 0);
  signal bram_addr_net: std_logic_vector(31 downto 0);
  signal bram_din_net: std_logic_vector(63 downto 0);
  signal bram_dout_net: std_logic_vector(63 downto 0);
  signal bram_en_net: std_logic;
  signal bram_reset_net: std_logic;
  signal bram_wen_net: std_logic_vector(7 downto 0);
  signal ce_1_sg_x98: std_logic;
  signal ce_8_sg_x3: std_logic;
  signal clk_1_sg_x98: std_logic;
  signal clk_8_sg_x3: std_logic;
  signal convert1_dout_net_x3: std_logic;
  signal convert2_dout_net_x5: std_logic_vector(8 downto 0);
  signal convert2_dout_net_x6: std_logic;
  signal convert6_dout_net_x3: std_logic_vector(1 downto 0);
  signal dac_tx_clk_net: std_logic;
  signal data_in_net: std_logic_vector(31 downto 0);
  signal data_in_x0_net: std_logic_vector(31 downto 0);
  signal data_in_x1_net: std_logic_vector(31 downto 0);
  signal data_in_x2_net: std_logic_vector(31 downto 0);
  signal data_in_x3_net: std_logic_vector(31 downto 0);
  signal data_in_x4_net: std_logic_vector(31 downto 0);
  signal data_in_x5_net: std_logic_vector(31 downto 0);
  signal data_out_net: std_logic_vector(31 downto 0);
  signal data_out_x0_net: std_logic_vector(31 downto 0);
  signal data_out_x1_net: std_logic_vector(31 downto 0);
  signal data_out_x2_net: std_logic_vector(31 downto 0);
  signal data_out_x3_net: std_logic_vector(31 downto 0);
  signal data_out_x4_net: std_logic_vector(31 downto 0);
  signal data_out_x5_net: std_logic_vector(31 downto 0);
  signal dbg_tx_running_net: std_logic;
  signal delay1_q_net_x2: std_logic;
  signal delay2_q_net_x1: std_logic;
  signal delay3_q_net_x7: std_logic;
  signal delay3_q_net_x8: std_logic;
  signal delay4_q_net_x1: std_logic;
  signal delay_q_net_x10: std_logic;
  signal delay_q_net_x11: std_logic;
  signal delay_q_net_x5: std_logic;
  signal dout_net: std_logic_vector(31 downto 0);
  signal dout_x0_net: std_logic_vector(31 downto 0);
  signal dout_x1_net: std_logic_vector(31 downto 0);
  signal dout_x2_net: std_logic_vector(31 downto 0);
  signal dout_x3_net: std_logic_vector(31 downto 0);
  signal dout_x4_net: std_logic_vector(31 downto 0);
  signal en_net: std_logic;
  signal en_x0_net: std_logic;
  signal en_x1_net: std_logic;
  signal en_x2_net: std_logic;
  signal en_x3_net: std_logic;
  signal en_x4_net: std_logic;
  signal en_x5_net: std_logic;
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4: std_logic_vector(15 downto 0);
  signal fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2: std_logic;
  signal fast_fourier_transform_8_0_s_axis_data_tready_net_x2: std_logic;
  signal fifo_dcount_net_x3: std_logic_vector(7 downto 0);
  signal logical1_y_net_x13: std_logic;
  signal logical1_y_net_x2: std_logic;
  signal logical1_y_net_x5: std_logic;
  signal logical2_y_net_x2: std_logic;
  signal logical_y_net_x3: std_logic;
  signal logical_y_net_x50: std_logic;
  signal logical_y_net_x7: std_logic;
  signal lsb_y_net_x1: std_logic;
  signal mux3_y_net_x1: std_logic_vector(11 downto 0);
  signal mux4_y_net_x1: std_logic_vector(11 downto 0);
  signal mux_y_net_x3: std_logic_vector(3 downto 0);
  signal mux_y_net_x7: std_logic;
  signal mux_y_net_x8: std_logic;
  signal phy_tx_done_net: std_logic;
  signal phy_tx_pkt_buf_net: std_logic_vector(3 downto 0);
  signal phy_tx_start_net: std_logic;
  signal phy_tx_started_net: std_logic;
  signal plb_ce_1_sg_x1: std_logic;
  signal plb_clk_1_sg_x1: std_logic;
  signal rc_phy_start_net: std_logic;
  signal rc_usr_rxen_net: std_logic;
  signal rc_usr_txen_net: std_logic;
  signal register2_q_net_x6: std_logic;
  signal register_q_net_x2: std_logic;
  signal reinterpret1_output_port_net_x2: std_logic_vector(15 downto 0);
  signal reinterpret2_output_port_net_x3: std_logic_vector(15 downto 0);
  signal reinterpret3_output_port_net_x3: std_logic_vector(15 downto 0);
  signal reinterpret_output_port_net_x2: std_logic_vector(15 downto 0);
  signal rfa_dac_i_net: std_logic_vector(11 downto 0);
  signal rfa_dac_q_net: std_logic_vector(11 downto 0);
  signal rfb_dac_i_net: std_logic_vector(11 downto 0);
  signal rfb_dac_q_net: std_logic_vector(11 downto 0);
  signal rx_sigs_invalid_net: std_logic;
  signal s_axi_araddr_net: std_logic_vector(31 downto 0);
  signal s_axi_arburst_net: std_logic_vector(1 downto 0);
  signal s_axi_arcache_net: std_logic_vector(3 downto 0);
  signal s_axi_arid_net: std_logic_vector(7 downto 0);
  signal s_axi_arlen_net: std_logic_vector(7 downto 0);
  signal s_axi_arlock_net: std_logic_vector(1 downto 0);
  signal s_axi_arprot_net: std_logic_vector(2 downto 0);
  signal s_axi_arready_net: std_logic;
  signal s_axi_arsize_net: std_logic_vector(2 downto 0);
  signal s_axi_arvalid_net: std_logic;
  signal s_axi_awaddr_net: std_logic_vector(31 downto 0);
  signal s_axi_awburst_net: std_logic_vector(1 downto 0);
  signal s_axi_awcache_net: std_logic_vector(3 downto 0);
  signal s_axi_awid_net: std_logic_vector(7 downto 0);
  signal s_axi_awlen_net: std_logic_vector(7 downto 0);
  signal s_axi_awlock_net: std_logic_vector(1 downto 0);
  signal s_axi_awprot_net: std_logic_vector(2 downto 0);
  signal s_axi_awready_net: std_logic;
  signal s_axi_awsize_net: std_logic_vector(2 downto 0);
  signal s_axi_awvalid_net: std_logic;
  signal s_axi_bid_net: std_logic_vector(7 downto 0);
  signal s_axi_bready_net: std_logic;
  signal s_axi_bresp_net: std_logic_vector(1 downto 0);
  signal s_axi_bvalid_net: std_logic;
  signal s_axi_rdata_net: std_logic_vector(31 downto 0);
  signal s_axi_rid_net: std_logic_vector(7 downto 0);
  signal s_axi_rlast_net: std_logic;
  signal s_axi_rready_net: std_logic;
  signal s_axi_rresp_net: std_logic_vector(1 downto 0);
  signal s_axi_rvalid_net: std_logic;
  signal s_axi_wdata_net: std_logic_vector(31 downto 0);
  signal s_axi_wlast_net: std_logic;
  signal s_axi_wready_net: std_logic;
  signal s_axi_wstrb_net: std_logic_vector(3 downto 0);
  signal s_axi_wvalid_net: std_logic;

begin
  axi_aresetn_net <= axi_aresetn;
  bram_din_net <= bram_din;
  ce_1_sg_x98 <= ce_1;
  ce_8_sg_x3 <= ce_8;
  clk_1_sg_x98 <= clk_1;
  clk_8_sg_x3 <= clk_8;
  dac_tx_clk_net <= dac_tx_clk;
  data_out_net <= data_out;
  data_out_x0_net <= data_out_x0;
  data_out_x1_net <= data_out_x1;
  data_out_x2_net <= data_out_x2;
  data_out_x3_net <= data_out_x3;
  data_out_x4_net <= data_out_x4;
  data_out_x5_net <= data_out_x5;
  dout_net <= dout;
  dout_x0_net <= dout_x0;
  dout_x1_net <= dout_x1;
  dout_x2_net <= dout_x2;
  dout_x3_net <= dout_x3;
  dout_x4_net <= dout_x4;
  phy_tx_pkt_buf_net <= phy_tx_pkt_buf;
  phy_tx_start_net <= phy_tx_start;
  plb_ce_1_sg_x1 <= plb_ce_1;
  plb_clk_1_sg_x1 <= plb_clk_1;
  rc_phy_start_net <= rc_phy_start;
  s_axi_araddr_net <= s_axi_araddr;
  s_axi_arburst_net <= s_axi_arburst;
  s_axi_arcache_net <= s_axi_arcache;
  s_axi_arid_net <= s_axi_arid;
  s_axi_arlen_net <= s_axi_arlen;
  s_axi_arlock_net <= s_axi_arlock;
  s_axi_arprot_net <= s_axi_arprot;
  s_axi_arsize_net <= s_axi_arsize;
  s_axi_arvalid_net <= s_axi_arvalid;
  s_axi_awaddr_net <= s_axi_awaddr;
  s_axi_awburst_net <= s_axi_awburst;
  s_axi_awcache_net <= s_axi_awcache;
  s_axi_awid_net <= s_axi_awid;
  s_axi_awlen_net <= s_axi_awlen;
  s_axi_awlock_net <= s_axi_awlock;
  s_axi_awprot_net <= s_axi_awprot;
  s_axi_awsize_net <= s_axi_awsize;
  s_axi_awvalid_net <= s_axi_awvalid;
  s_axi_bready_net <= s_axi_bready;
  s_axi_rready_net <= s_axi_rready;
  s_axi_wdata_net <= s_axi_wdata;
  s_axi_wlast_net <= s_axi_wlast;
  s_axi_wstrb_net <= s_axi_wstrb;
  s_axi_wvalid_net <= s_axi_wvalid;
  bram_addr <= bram_addr_net;
  bram_dout <= bram_dout_net;
  bram_en <= bram_en_net;
  bram_reset <= bram_reset_net;
  bram_wen <= bram_wen_net;
  data_in <= data_in_net;
  data_in_x0 <= data_in_x0_net;
  data_in_x1 <= data_in_x1_net;
  data_in_x2 <= data_in_x2_net;
  data_in_x3 <= data_in_x3_net;
  data_in_x4 <= data_in_x4_net;
  data_in_x5 <= data_in_x5_net;
  dbg_tx_running <= dbg_tx_running_net;
  en <= en_net;
  en_x0 <= en_x0_net;
  en_x1 <= en_x1_net;
  en_x2 <= en_x2_net;
  en_x3 <= en_x3_net;
  en_x4 <= en_x4_net;
  en_x5 <= en_x5_net;
  phy_tx_done <= phy_tx_done_net;
  phy_tx_started <= phy_tx_started_net;
  rc_usr_rxen <= rc_usr_rxen_net;
  rc_usr_txen <= rc_usr_txen_net;
  rfa_dac_i <= rfa_dac_i_net;
  rfa_dac_q <= rfa_dac_q_net;
  rfb_dac_i <= rfb_dac_i_net;
  rfb_dac_q <= rfb_dac_q_net;
  rx_sigs_invalid <= rx_sigs_invalid_net;
  s_axi_arready <= s_axi_arready_net;
  s_axi_awready <= s_axi_awready_net;
  s_axi_bid <= s_axi_bid_net;
  s_axi_bresp <= s_axi_bresp_net;
  s_axi_bvalid <= s_axi_bvalid_net;
  s_axi_rdata <= s_axi_rdata_net;
  s_axi_rid <= s_axi_rid_net;
  s_axi_rlast <= s_axi_rlast_net;
  s_axi_rresp <= s_axi_rresp_net;
  s_axi_rvalid <= s_axi_rvalid_net;
  s_axi_wready <= s_axi_wready_net;

  bit_source_8a38dc99ff: entity work.bit_source_entity_8a38dc99ff
    port map (
      b_15_8 => b_15_8_y_net_x3,
      b_23_16 => b_23_16_y_net_x2,
      b_7_0 => b_7_0_y_net_x4,
      bram_din => bram_din_net,
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      convert2 => convert2_dout_net_x6,
      done => delay3_q_net_x8,
      fifo => fifo_dcount_net_x3,
      mux => mux_y_net_x3,
      tx_reset => logical_y_net_x50,
      tx_start => logical_y_net_x7,
      addr_gen => delay3_q_net_x7,
      bit => mux_y_net_x7,
      bit_valid => delay_q_net_x5,
      bram_if_64b => bram_addr_net,
      bram_if_64b_x0 => bram_en_net,
      bram_if_64b_x1 => bram_reset_net,
      bram_if_64b_x2 => bram_dout_net,
      bram_if_64b_x3 => bram_wen_net,
      data_pad_fcs => logical1_y_net_x5,
      signal_capture => convert2_dout_net_x5,
      signal_capture_x0 => convert6_dout_net_x3,
      signal_capture_x1 => b_2_1_y_net_x1,
      signal_decode_error => register_q_net_x2,
      tail => delay4_q_net_x1
    );

  edk_processor_de00edcbbe: entity work.edk_processor_entity_de00edcbbe
    port map (
      axi_aresetn => axi_aresetn_net,
      from_register => data_out_net,
      plb_ce_1 => plb_ce_1_sg_x1,
      plb_clk_1 => plb_clk_1_sg_x1,
      s_axi_araddr => s_axi_araddr_net,
      s_axi_arburst => s_axi_arburst_net,
      s_axi_arcache => s_axi_arcache_net,
      s_axi_arid => s_axi_arid_net,
      s_axi_arlen => s_axi_arlen_net,
      s_axi_arlock => s_axi_arlock_net,
      s_axi_arprot => s_axi_arprot_net,
      s_axi_arsize => s_axi_arsize_net,
      s_axi_arvalid => s_axi_arvalid_net,
      s_axi_awaddr => s_axi_awaddr_net,
      s_axi_awburst => s_axi_awburst_net,
      s_axi_awcache => s_axi_awcache_net,
      s_axi_awid => s_axi_awid_net,
      s_axi_awlen => s_axi_awlen_net,
      s_axi_awlock => s_axi_awlock_net,
      s_axi_awprot => s_axi_awprot_net,
      s_axi_awsize => s_axi_awsize_net,
      s_axi_awvalid => s_axi_awvalid_net,
      s_axi_bready => s_axi_bready_net,
      s_axi_rready => s_axi_rready_net,
      s_axi_wdata => s_axi_wdata_net,
      s_axi_wlast => s_axi_wlast_net,
      s_axi_wstrb => s_axi_wstrb_net,
      s_axi_wvalid => s_axi_wvalid_net,
      to_register => dout_net,
      to_register1 => dout_x0_net,
      to_register2 => dout_x1_net,
      to_register3 => dout_x2_net,
      to_register4 => dout_x3_net,
      to_register5 => dout_x4_net,
      memmap_x0 => s_axi_arready_net,
      memmap_x1 => s_axi_awready_net,
      memmap_x10 => s_axi_wready_net,
      memmap_x11 => data_in_net,
      memmap_x12 => en_net,
      memmap_x13 => data_in_x0_net,
      memmap_x14 => en_x0_net,
      memmap_x15 => data_in_x1_net,
      memmap_x16 => en_x1_net,
      memmap_x17 => data_in_x2_net,
      memmap_x18 => en_x2_net,
      memmap_x19 => data_in_x3_net,
      memmap_x2 => s_axi_bid_net,
      memmap_x20 => en_x3_net,
      memmap_x21 => data_in_x4_net,
      memmap_x22 => en_x4_net,
      memmap_x3 => s_axi_bresp_net,
      memmap_x4 => s_axi_bvalid_net,
      memmap_x5 => s_axi_rdata_net,
      memmap_x6 => s_axi_rid_net,
      memmap_x7 => s_axi_rlast_net,
      memmap_x8 => s_axi_rresp_net,
      memmap_x9 => s_axi_rvalid_net
    );

  fft_b2c6e5af27: entity work.fft_entity_b2c6e5af27
    port map (
      b_15_8 => b_15_8_y_net_x3,
      b_29_24 => b_29_24_y_net_x1,
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      data_in_tlast => logical2_y_net_x2,
      data_in_tvalid => axi_fifo_m_axis_tvalid_net_x2,
      i_in => reinterpret2_output_port_net_x3,
      last_sym => logical1_y_net_x2,
      q_in => reinterpret3_output_port_net_x3,
      tx_reset => logical_y_net_x50,
      data_in_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x2,
      data_out_tvalid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2,
      i_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4,
      last_sym_x0 => logical_y_net_x3,
      q_out => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4
    );

  fifo_c992f1a4af: entity work.fifo_entity_c992f1a4af
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      data_tvalid => delay_q_net_x10,
      fft_tready => fast_fourier_transform_8_0_s_axis_data_tready_net_x2,
      i => mux3_y_net_x1,
      last_samp => delay1_q_net_x2,
      last_sym => delay3_q_net_x8,
      q => mux4_y_net_x1,
      tx_reset => logical_y_net_x50,
      fft_tdata_im => reinterpret3_output_port_net_x3,
      fft_tdata_re => reinterpret2_output_port_net_x3,
      fft_tlast => logical2_y_net_x2,
      fft_tvalid => axi_fifo_m_axis_tvalid_net_x2,
      fifo_tready => axi_fifo_s_axis_tready_net_x2,
      last_sym_x0 => logical1_y_net_x2
    );

  interleave_modulate_1e78258d30: entity work.\interleave___modulate_entity_1e78258d30\
    port map (
      b_7_0 => b_7_0_y_net_x4,
      bit => mux_y_net_x8,
      bit_source => delay3_q_net_x7,
      bit_source_x0 => convert2_dout_net_x5,
      bit_valid => delay_q_net_x11,
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      fifo_in_ready => axi_fifo_s_axis_tready_net_x2,
      logical => logical_y_net_x50,
      signal_mod_sel => b_2_1_y_net_x1,
      last_sym => delay3_q_net_x8,
      x_i => mux3_y_net_x1,
      x_iq_last => delay1_q_net_x2,
      x_iq_valid => delay_q_net_x10,
      x_q => mux4_y_net_x1
    );

  preamble_outputs_82fcc722dc: entity work.\preamble___outputs_entity_82fcc722dc\
    port map (
      b_2 => b_2_y_net_x1,
      b_3 => b_3_y_net_x1,
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      fft_i => fast_fourier_transform_8_0_m_axis_data_tdata_xk_re_net_x4,
      fft_i_q_valid => fast_fourier_transform_8_0_m_axis_data_tvalid_net_x2,
      fft_q => fast_fourier_transform_8_0_m_axis_data_tdata_xk_im_net_x4,
      last_sym => logical_y_net_x3,
      reinterpret => reinterpret_output_port_net_x2,
      reinterpret1 => reinterpret1_output_port_net_x2,
      tx_iq_samp_ce => convert2_dout_net_x6,
      tx_reset => logical_y_net_x50,
      tx_start => logical_y_net_x7,
      dac_outputs => rfa_dac_i_net,
      dac_outputs_x0 => rfa_dac_q_net,
      dac_outputs_x1 => rfb_dac_i_net,
      dac_outputs_x2 => rfb_dac_q_net,
      last_samp_output_to_dacs => delay2_q_net_x1,
      output_fifo_occ => fifo_dcount_net_x3
    );

  registers_2d8965b1e5: entity work.registers_entity_2d8965b1e5
    port map (
      from_register1 => data_out_x0_net,
      from_register2 => data_out_x1_net,
      from_register3 => data_out_x2_net,
      from_register4 => data_out_x3_net,
      from_register5 => data_out_x4_net,
      from_register6 => data_out_x5_net,
      register2 => register2_q_net_x6,
      constant_x1 => en_x5_net,
      regtx_anta_tx_en => b_2_y_net_x1,
      regtx_antb_tx_en => b_3_y_net_x1,
      regtx_cp_len => b_15_8_y_net_x3,
      regtx_fft_scaling => b_29_24_y_net_x1,
      regtx_num_sc => b_7_0_y_net_x4,
      regtx_pkt_buf_addr_offset => b_23_16_y_net_x2,
      regtx_pkt_buf_sel => b_3_0_y_net_x1,
      regtx_posttx_extension => b_7_0_1_y_net_x2,
      regtx_posttx_rf_en_extension => b_15_8_1_y_net_x2,
      regtx_posttx_rxsig_valid => b_23_16_y_net_x1,
      regtx_rc_rxen_enable => b_0_1_y_net_x1,
      regtx_reset => b_31_y_net_x0,
      regtx_reset_scrambling_lfsr_perpkt => b_1_y_net_x2,
      regtx_scaling_payload => reinterpret1_output_port_net_x2,
      regtx_scaling_preamble => reinterpret_output_port_net_x2,
      regtx_start_direct => lsb_y_net_x1,
      regtx_start_indirect => b_1_y_net_x3,
      status_bits => data_in_x5_net
    );

  resets_24d0a1b807: entity work.resets_entity_24d0a1b807
    port map (
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      last_samp_output_to_dacs => delay2_q_net_x1,
      regtx_reset => b_31_y_net_x0,
      signal_decode_error => register_q_net_x2,
      tx_force_reset => convert1_dout_net_x3,
      tx_phy_done => logical1_y_net_x13,
      tx_reset => logical_y_net_x50
    );

  scramble_encode_5f70e14e46: entity work.\scramble___encode_entity_5f70e14e46\
    port map (
      bit => mux_y_net_x7,
      bit_source => convert6_dout_net_x3,
      bit_valid => delay_q_net_x5,
      ce_1 => ce_1_sg_x98,
      clk_1 => clk_1_sg_x98,
      data_pad_fcs => logical1_y_net_x5,
      registers => b_1_y_net_x2,
      tail => delay4_q_net_x1,
      tx_reset => logical_y_net_x50,
      enc_bit => mux_y_net_x8,
      enc_bit_valid => delay_q_net_x11
    );

  start_ctrl_3ba2a032ad: entity work.start_ctrl_entity_3ba2a032ad
    port map (
      ce_1 => ce_1_sg_x98,
      ce_8 => ce_8_sg_x3,
      clk_1 => clk_1_sg_x98,
      clk_8 => clk_8_sg_x3,
      dac_tx_clk => dac_tx_clk_net,
      phy_tx_pkt_buf => phy_tx_pkt_buf_net,
      phy_tx_start => phy_tx_start_net,
      rc_phy_start => rc_phy_start_net,
      registers => b_15_8_1_y_net_x2,
      registers_x0 => b_23_16_y_net_x1,
      registers_x1 => b_3_0_y_net_x1,
      registers_x2 => b_7_0_1_y_net_x2,
      regtx_rc_rxen_enable => b_0_1_y_net_x1,
      regtx_start_direct => lsb_y_net_x1,
      regtx_start_indirect => b_1_y_net_x3,
      tx_force_reset => convert1_dout_net_x3,
      tx_phy_done => logical1_y_net_x13,
      negedge_x0 => phy_tx_done_net,
      phy_start => logical_y_net_x7,
      posedge2 => phy_tx_started_net,
      register1_x0 => dbg_tx_running_net,
      register2_x0 => rx_sigs_invalid_net,
      register4_x0 => rc_usr_rxen_net,
      register5_x0 => rc_usr_txen_net,
      regtx_tx_running => register2_q_net_x6,
      tx_iq_samp_ce => convert2_dout_net_x6,
      tx_pkt_buf_sel => mux_y_net_x3
    );

end structural;
